module Loading_Screen (
    input logic CLK, RESET, Loading_Text,
    input logic [9:0] DrawX, DrawY,
    output logic loading_active
);



//logic zeroidx, oneidx, twoidx, threeidx, fouridx, fiveidx, sixidx, sevenidx, eightidx, nineidx, tenidx, elevenidx;
//logic twelveidx, thirteenidx, fourteenidx, fifteenidx, sixteenidx, seventeenidx, eighteenidx, nineteenidx;
logic [9:0] mod8;
assign mod8 = (DrawY + 8) % 16;


always_comb begin : print_letters 
    
    
    if(Loading_Text) begin
        if( (292 > DrawX) & (DrawX >= 284) & (376 > DrawY) & (DrawY>= 360) ) begin
            logic [9:0] bah;
            bah = DrawX-284;

            loading_active = LetterL[mod8[3:0]][bah[2:0]];
            
        end

        else if( (300 > DrawX) & (DrawX >= 292) & (376 > DrawY) & (DrawY>= 360) ) begin
            logic [9:0] bah;
            bah = DrawX-292;

            loading_active = LetterO[mod8[3:0]][bah[2:0]];
            
        end   

        else if( (308 > DrawX) & (DrawX >= 300) & (376 > DrawY) & (DrawY>= 360) ) begin
            logic [9:0] bah;
            bah = DrawX-300;

            loading_active = LetterA[mod8[3:0]][bah[2:0]];
            
        end

        else if( (316 > DrawX) & (DrawX >= 308) & (376 > DrawY) & (DrawY>= 360) ) begin
            logic [9:0] bah;
            bah = DrawX-308;

            loading_active = LetterD[mod8[3:0]][bah[2:0]];
            
        end  

        else if( (324 > DrawX) & (DrawX >= 316) & (376 > DrawY) & (DrawY>= 360) ) begin
            logic [9:0] bah;
            bah = DrawX-316;

            loading_active = LetterI[mod8[3:0]][bah[2:0]];
            
        end 

        else if( (332 > DrawX) & (DrawX >= 324) & (376 > DrawY) & (DrawY>= 360) ) begin
            logic [9:0] bah;
            bah = DrawX-324;

            loading_active = LetterN[mod8[3:0]][bah[2:0]];
            
        end 

        else if( (340 > DrawX) & (DrawX >= 332) & (376 > DrawY) & (DrawY>= 360) ) begin
            logic [9:0] bah;
            bah = DrawX-332;

            loading_active = LetterG[mod8[3:0]][bah[2:0]];
            
        end 

        else if( (348 > DrawX) & (DrawX >= 340) & (376 > DrawY) & (DrawY>= 360) ) begin
            logic [9:0] bah;
            bah = DrawX-340;

            loading_active = LetterPeriod[mod8[3:0]][bah[2:0]];
            
        end 
        
        else if( (356 > DrawX) & (DrawX >= 348) & (376 > DrawY) & (DrawY>= 360) ) begin
            logic [9:0] bah;
            bah = DrawX-326;

            loading_active = LetterPeriod[mod8[3:0]][bah[2:0]];
            
        end 

        else if( (364 > DrawX) & (DrawX >= 356) & (376 > DrawY) & (DrawY>= 360) ) begin
            logic [9:0] bah;
            bah = DrawX-356;

            loading_active = LetterPeriod[mod8[3:0]][bah[2:0]];
            
        end   
        else
            loading_active = 0; 

    end
    else begin
        loading_active = 0;
    end
    
end


    parameter bit LetterN[16][8] = '{
        '{0,0,0,0,0,0,0,0}, // 0
        '{0,0,0,0,0,0,0,0}, // 1
        '{1,1,0,0,0,1,1,0}, // 2 **   **
        '{1,1,1,0,0,1,1,0}, // 3 ***  **
        '{1,1,1,1,0,1,1,0}, // 4 **** **
        '{1,1,1,1,1,1,1,0}, // 5 *******
        '{1,1,0,1,1,1,1,0}, // 6 ** ****
        '{1,1,0,0,1,1,1,0}, // 7 **  ***
        '{1,1,0,0,0,1,1,0}, // 8 **   **
        '{1,1,0,0,0,1,1,0}, // 9 **   **
        '{1,1,0,0,0,1,1,0}, // a **   **
        '{1,1,0,0,0,1,1,0}, // b **   **
        '{0,0,0,0,0,0,0,0}, // c
        '{0,0,0,0,0,0,0,0}, // d
        '{0,0,0,0,0,0,0,0}, // e
        '{0,0,0,0,0,0,0,0} // f
    };
    

    parameter bit LetterO[16][8] = '{
        '{0,0,0,0,0,0,0,0}, // 0
        '{0,0,0,0,0,0,0,0}, // 1
        '{0,1,1,1,1,1,0,0}, // 2  *****
        '{1,1,0,0,0,1,1,0}, // 3 **   **
        '{1,1,0,0,0,1,1,0}, // 4 **   **
        '{1,1,0,0,0,1,1,0}, // 5 **   **
        '{1,1,0,0,0,1,1,0}, // 6 **   **
        '{1,1,0,0,0,1,1,0}, // 7 **   **
        '{1,1,0,0,0,1,1,0}, // 8 **   **
        '{1,1,0,0,0,1,1,0}, // 9 **   **
        '{1,1,0,0,0,1,1,0}, // a **   **
        '{0,1,1,1,1,1,0,0}, // b  *****
        '{0,0,0,0,0,0,0,0}, // c
        '{0,0,0,0,0,0,0,0}, // d
        '{0,0,0,0,0,0,0,0}, // e
        '{0,0,0,0,0,0,0,0} // f
    };
    parameter bit LetterA[16][8] = '{
        '{0,0,0,0,0,0,0,0}, // 0
        '{0,0,0,0,0,0,0,0}, // 1
        '{0,0,0,1,0,0,0,0}, // 2    *
        '{0,0,1,1,1,0,0,0}, // 3   ***
        '{0,1,1,0,1,1,0,0}, // 4  ** **
        '{1,1,0,0,0,1,1,0}, // 5 **   **
        '{1,1,0,0,0,1,1,0}, // 6 **   **
        '{1,1,1,1,1,1,1,0}, // 7 *******
        '{1,1,0,0,0,1,1,0}, // 8 **   **
        '{1,1,0,0,0,1,1,0}, // 9 **   **
        '{1,1,0,0,0,1,1,0}, // a **   **
        '{1,1,0,0,0,1,1,0}, // b **   **
        '{0,0,0,0,0,0,0,0}, // c
        '{0,0,0,0,0,0,0,0}, // d
        '{0,0,0,0,0,0,0,0}, // e
        '{0,0,0,0,0,0,0,0} // f
    };
    parameter bit LetterG[16][8] = '{
        '{0,0,0,0,0,0,0,0}, // 0
        '{0,0,0,0,0,0,0,0}, // 1
        '{0,0,1,1,1,1,0,0}, // 2   ****
        '{0,1,1,0,0,1,1,0}, // 3  **  **
        '{1,1,0,0,0,0,1,0}, // 4 **    *
        '{1,1,0,0,0,0,0,0}, // 5 **
        '{1,1,0,0,0,0,0,0}, // 6 **
        '{1,1,0,1,1,1,1,0}, // 7 ** ****
        '{1,1,0,0,0,1,1,0}, // 8 **   **
        '{1,1,0,0,0,1,1,0}, // 9 **   **
        '{0,1,1,0,0,1,1,0}, // a  **  **
        '{0,0,1,1,1,0,1,0}, // b   *** *
        '{0,0,0,0,0,0,0,0}, // c
        '{0,0,0,0,0,0,0,0}, // d
        '{0,0,0,0,0,0,0,0}, // e
        '{0,0,0,0,0,0,0,0} // f
    };
    parameter bit LetterL[16][8] = '{
        '{0,0,0,0,0,0,0,0}, // 0
        '{0,0,0,0,0,0,0,0}, // 1
        '{1,1,1,1,0,0,0,0}, // 2 ****
        '{0,1,1,0,0,0,0,0}, // 3  **
        '{0,1,1,0,0,0,0,0}, // 4  **
        '{0,1,1,0,0,0,0,0}, // 5  **
        '{0,1,1,0,0,0,0,0}, // 6  **
        '{0,1,1,0,0,0,0,0}, // 7  **
        '{0,1,1,0,0,0,0,0}, // 8  **
        '{0,1,1,0,0,0,1,0}, // 9  **   *
        '{0,1,1,0,0,1,1,0}, // a  **  **
        '{1,1,1,1,1,1,1,0}, // b *******
        '{0,0,0,0,0,0,0,0}, // c
        '{0,0,0,0,0,0,0,0}, // d
        '{0,0,0,0,0,0,0,0}, // e
        '{0,0,0,0,0,0,0,0} // f
    };
    parameter bit LetterD[16][8] = '{
        '{0,0,0,0,0,0,0,0}, // 0
        '{0,0,0,0,0,0,0,0}, // 1
        '{1,1,1,1,1,0,0,0}, // 2 *****
        '{0,1,1,0,1,1,0,0}, // 3  ** **
        '{0,1,1,0,0,1,1,0}, // 4  **  **
        '{0,1,1,0,0,1,1,0}, // 5  **  **
        '{0,1,1,0,0,1,1,0}, // 6  **  **
        '{0,1,1,0,0,1,1,0}, // 7  **  **
        '{0,1,1,0,0,1,1,0}, // 8  **  **
        '{0,1,1,0,0,1,1,0}, // 9  **  **
        '{0,1,1,0,1,1,0,0}, // a  ** **
        '{1,1,1,1,1,0,0,0}, // b *****
        '{0,0,0,0,0,0,0,0}, // c
        '{0,0,0,0,0,0,0,0}, // d
        '{0,0,0,0,0,0,0,0}, // e
        '{0,0,0,0,0,0,0,0} // f
    };
    parameter bit LetterI[16][8] = '{
        '{0,0,0,0,0,0,0,0}, // 0
        '{0,0,0,0,0,0,0,0}, // 1
        '{0,0,1,1,1,1,0,0}, // 2   ****
        '{0,0,0,1,1,0,0,0}, // 3    **
        '{0,0,0,1,1,0,0,0}, // 4    **
        '{0,0,0,1,1,0,0,0}, // 5    **
        '{0,0,0,1,1,0,0,0}, // 6    **
        '{0,0,0,1,1,0,0,0}, // 7    **
        '{0,0,0,1,1,0,0,0}, // 8    **
        '{0,0,0,1,1,0,0,0}, // 9    **
        '{0,0,0,1,1,0,0,0}, // a    **
        '{0,0,1,1,1,1,0,0}, // b   ****
        '{0,0,0,0,0,0,0,0}, // c
        '{0,0,0,0,0,0,0,0}, // d
        '{0,0,0,0,0,0,0,0}, // e
        '{0,0,0,0,0,0,0,0}// f
    };
    parameter bit LetterPeriod[16][8] = '{
        '{0,0,0,0,0,0,0,0}, // 0
        '{0,0,0,0,0,0,0,0}, // 1
        '{0,0,0,0,0,0,0,0}, // 2
        '{0,0,0,0,0,0,0,0}, // 3
        '{0,0,0,0,0,0,0,0}, // 4
        '{0,0,0,0,0,0,0,0}, // 5
        '{0,0,0,0,0,0,0,0}, // 6
        '{0,0,0,0,0,0,0,0}, // 7
        '{0,0,0,0,0,0,0,0}, // 8
        '{0,0,0,0,0,0,0,0}, // 9
        '{0,0,0,1,1,0,0,0}, // a    **
        '{0,0,0,1,1,0,0,0}, // b    **
        '{0,0,0,0,0,0,0,0}, // c
        '{0,0,0,0,0,0,0,0}, // d
        '{0,0,0,0,0,0,0,0}, // e
        '{0,0,0,0,0,0,0,0} // f
    };
     

endmodule