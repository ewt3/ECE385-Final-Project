module Jerry(
input CLK,
input logic RESET, Pause, invincibility,
input logic frame_clk, switch, dead,
input logic [7:0] KeyCodes,
input logic [9:0] DrawX, DrawY, 
output logic active, offscreen,
output logic [11:0] Color,
output logic [9:0] JerryX, JerryY  //, JerrywidthEnd, JerryheightEnd
);


//local variables
logic [9:0] Jerry_X_Pos, Jerry_X_Motion, Jerry_Y_Pos, Jerry_Y_Motion, width, height, widthEnd, heightEnd;
//logic [8:0] movement_counter;
	
parameter [9:0] Jerry_X_Center=320;  // Center position on the X axis
parameter [9:0] Jerry_Y_Center=240;  // Center position on the Y axis
parameter [9:0] Jerry_X_Min=0;       // Leftmost point on the X axis
parameter [9:0] Jerry_X_Max=639;     // Rightmost point on the X axis
parameter [9:0] Jerry_Y_Min=0;       // Topmost point on the Y axis
parameter [9:0] Jerry_Y_Max=479;     // Bottommost point on the Y axis
logic [9:0] Jerry_X_Step;     // Step size on the X axis
logic [9:0] Jerry_Y_Step;      // Step size on the Y axis

always_comb begin
	if(invincibility) begin
		Jerry_X_Step = 10;
		Jerry_Y_Step = 10;
	end
	else begin
		Jerry_X_Step = 3;
		Jerry_Y_Step = 3;
	end

end


assign width = 25;
assign height = 35;

assign JerryX = Jerry_X_Pos;
assign JerryY = Jerry_Y_Pos;



always_comb begin : Active_Logic // can be simplified at expense of readibility
	widthEnd = width + Jerry_X_Pos;
	heightEnd = height + Jerry_Y_Pos;
	if(dead) begin
		if(deadCounter[25])begin
			if(	(DrawX >= Jerry_X_Pos) & (DrawX < Jerry_X_Pos + 37) & 
			(DrawY >= Jerry_Y_Pos) & (DrawY < Jerry_Y_Pos + 29) ) begin
				if((Color == 12'h111))
					active = 0;
				else	
					active = 1;
			end 
			else begin
				active = 0;
			end
		end else begin
			if(	(DrawX >= Jerry_X_Pos) & (DrawX < Jerry_X_Pos + 29) & 
			(DrawY >= Jerry_Y_Pos) & (DrawY < Jerry_Y_Pos + 37) ) begin
				if((Color == 12'h111))
					active = 0;
				else	
					active = 1;
			end 
			else begin
				active = 0;
			end
		end
	end
	else begin
		if(	(DrawX >= Jerry_X_Pos) & (DrawX < widthEnd) & 
			(DrawY >= Jerry_Y_Pos) & (DrawY < heightEnd) ) begin
				if((Color == 12'h111))
					active = 0;
				else	
					active = 1;
			end 
		else begin
			active = 0;
		end
	end
		
end






logic [25:0] deadCounter;
always_ff @( posedge CLK or posedge RESET) begin : AnimationCounter
	if(RESET)begin
		deadCounter <= 0;
	end else begin
		if(dead)
			if(deadCounter[25])
				deadCounter <= deadCounter;
			else
				deadCounter <= deadCounter + 1;
		else
			deadCounter <= 0;
	end
end

logic [6:0] indx, indy;
always_comb begin : Pallete_Assignment
	indx = DrawX - Jerry_X_Pos;
	indy = DrawY - Jerry_Y_Pos;
	if(dead) begin
		if(deadCounter[25])
			Color = DeadJerryColors1[indy][indx];
		else
			Color = DeadJerryColors2[indy][indx];
	end else begin
		if(switch)
			//pallete = JerryColors1[indy][indx];
			Color = JerryColors1[indy][indx];
		else
			//pallete = JerryColors2[indy][indx];
			Color = JerryColors2[indy][indx];
	end
end






//Jerry definition
parameter bit [11:0] JerryColors1 [35][25] = '{
'{273,273,273,0,0,0,273,273,273,273,273,273,273,273,273,0,0,0,0,0,0,0,273,273,273},
'{273,273,0,0,2403,0,0,273,273,273,273,273,273,273,0,0,2403,2403,2403,2403,2403,0,0,273,273},
'{273,273,0,2403,2403,2403,0,273,273,273,273,273,273,0,0,2403,2403,4005,4005,4005,4005,2403,0,0,273},
'{273,273,0,2403,2403,2403,0,0,0,0,0,0,0,0,2403,2403,0,4005,4005,4005,4005,4005,2403,0,0},
'{273,273,0,2403,2403,0,0,2403,2403,2403,2403,2403,2403,0,0,2403,0,4005,4005,4005,4005,4005,4005,2403,0},
'{273,273,0,2403,2403,0,2403,2403,2403,2403,2403,2403,2403,2403,0,2403,0,0,4005,4005,4005,4005,4005,2403,0},
'{273,273,0,0,0,0,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,0,0,4005,4005,4005,2403,2403,0},
'{273,273,273,0,0,2131,0,0,2403,2403,2403,0,0,2403,2403,2403,2403,2403,0,0,0,2403,2403,0,0},
'{273,273,273,273,0,2403,0,0,2403,2403,2403,0,0,2403,2403,2403,2403,2403,2403,2403,2403,2403,0,0,273},
'{0,0,273,0,0,2403,0,0,2403,2403,2403,0,0,2403,2403,2403,2403,2403,2403,2403,0,0,0,273,273},
'{3549,0,0,0,0,2403,2403,2403,2403,2403,2403,2403,2403,0,0,0,0,0,2403,2403,0,273,273,273,273},
'{273,273,273,0,4005,4005,0,0,0,4005,4005,0,0,0,2403,2403,2403,2403,2403,2403,0,273,273,273,273},
'{273,0,0,0,0,4005,4005,4005,4005,4005,4005,4005,2403,2403,2403,2403,2403,2403,2403,2403,0,273,273,273,273},
'{0,0,273,0,4005,4005,0,4005,4005,0,4005,0,0,0,0,2403,2403,2403,2403,2403,0,273,273,273,273},
'{0,273,273,0,0,4005,4005,0,0,4005,4005,4005,4005,4005,0,0,2403,2403,2403,2403,0,273,273,273,273},
'{273,273,273,273,0,0,0,4005,4005,4005,4005,4005,4005,4005,2403,2403,2403,0,2403,2403,0,0,273,273,273},
'{273,273,273,273,273,273,0,0,0,4005,4005,4005,4005,2403,2403,0,0,0,2403,2403,2403,0,273,273,273},
'{273,273,273,273,0,0,0,2403,0,0,0,0,0,0,0,0,2403,2403,2403,2403,2403,0,0,273,273},
'{273,273,273,0,0,0,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,0,0,273},
'{273,273,0,0,2403,0,2403,2403,4005,4005,2403,2403,4005,4005,4005,2403,2403,2403,2403,2403,2403,2403,2403,0,273},
'{273,0,0,2403,2403,0,2403,4005,4005,4005,4005,4005,4005,4005,4005,2403,2403,2403,2403,2403,2403,2403,2403,0,0},
'{0,0,2403,2403,2403,0,2403,4005,4005,4005,4005,4005,4005,4005,4005,4005,2403,2403,2403,2403,2403,2403,2403,2403,0},
'{0,0,2403,2403,2403,0,2403,4005,4005,4005,4005,4005,4005,4005,4005,4005,4005,2403,2403,2403,0,2403,2403,2403,0},
'{273,0,0,2403,2403,0,2403,4005,4005,4005,4005,4005,4005,4005,4005,4005,4005,2403,2403,2403,0,0,2403,2403,0},
'{273,273,0,0,0,0,2403,4005,4005,4005,4005,4005,4005,4005,4005,4005,4005,2403,2403,2403,0,0,0,0,0},
'{273,273,273,273,273,0,2403,4005,4005,4005,4005,4005,4005,4005,4005,4005,4005,2403,2403,2403,0,273,273,273,273},
'{273,273,273,273,273,0,0,4005,4005,4005,4005,4005,4005,4005,4005,4005,4005,2403,2403,2403,0,273,273,273,273},
'{273,273,273,273,273,0,0,0,4005,4005,4005,4005,4005,4005,4005,4005,2403,2403,2403,2403,0,273,273,273,273},
'{273,273,273,273,273,0,2403,0,0,0,4005,4005,4005,4005,2403,2403,2403,2403,2403,2403,0,0,273,273,273},
'{273,273,273,273,273,0,2403,2403,2403,0,0,0,0,0,2403,2403,2403,2403,2403,2403,0,0,0,273,273},
'{273,273,273,273,273,0,2403,2403,2403,2403,2403,0,273,0,2403,2403,2403,2403,2403,2403,0,273,0,0,0},
'{273,273,273,273,273,0,0,2403,2403,2403,2403,0,273,0,2403,2403,2403,2403,2403,0,0,273,273,273,273},
'{273,273,273,273,273,273,0,2403,2403,2403,0,0,273,273,0,2403,2403,2403,2403,0,273,273,273,273,273},
'{273,273,273,273,273,273,0,0,2403,2403,0,273,273,273,0,0,2403,2403,0,0,273,273,273,273,273},
'{273,273,273,273,273,273,273,0,0,0,0,273,273,273,273,273,0,0,0,273,273,273,273,273,273}
};



parameter bit [11:0] JerryColors2 [35][25] = '{
'{273,273,273,0,0,0,273,273,273,273,273,273,273,273,273,0,0,0,0,0,0,0,273,273,273},
'{273,273,0,0,2403,0,0,273,273,273,273,273,273,273,0,0,2403,2403,2403,2403,2403,0,0,273,273},
'{273,273,0,2403,2403,2403,0,273,273,273,273,273,273,0,0,2403,2403,4005,4005,4005,4005,2403,0,0,273},
'{273,273,0,2403,2403,2403,0,0,0,0,0,0,0,0,2403,2403,0,4005,4005,4005,4005,4005,2403,0,0},
'{273,273,0,2403,2403,0,0,2403,2403,2403,2403,2403,2403,0,0,2403,0,4005,4005,4005,4005,4005,4005,2403,0},
'{273,273,0,2403,2403,0,2403,2403,2403,2403,2403,2403,2403,2403,0,2403,0,0,4005,4005,4005,4005,4005,2403,0},
'{273,273,0,0,0,0,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,0,0,4005,4005,4005,2403,2403,0},
'{273,273,273,0,0,2403,0,0,2403,2403,2403,0,0,2403,2403,2403,2403,2403,0,0,0,2403,2403,0,0},
'{273,273,273,273,0,2403,0,0,2403,2403,2403,0,0,2403,2403,2403,2403,2403,2403,2403,2403,2403,0,0,273},
'{273,273,273,0,0,2403,0,0,2403,2403,2403,0,0,2403,2403,2403,2403,2403,2403,2403,0,0,0,273,273},
'{0,0,0,0,0,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,0,273,273,273,273},
'{273,273,273,0,4005,4005,0,0,0,4005,4005,0,0,0,0,0,0,2403,2403,2403,0,273,273,273,273},
'{273,0,0,0,0,4005,4005,4005,4005,4005,4005,4005,2403,2403,2403,2403,2403,2403,2403,2403,0,273,273,273,273},
'{0,0,0,0,4005,4005,0,4005,4005,0,4005,0,0,0,2403,2403,2403,2403,2403,2403,0,273,273,273,273},
'{0,273,273,0,0,4005,4005,0,0,4005,4005,4005,4005,0,0,2403,2403,2403,2403,2403,0,273,273,273,273},
'{273,273,273,273,0,0,0,4005,4005,4005,4005,4005,4005,4005,0,2403,2403,0,2403,2403,0,0,273,273,273},
'{273,273,273,273,273,273,0,0,0,4005,4005,4005,4005,2403,2403,0,0,0,2403,2403,2403,0,273,273,273},
'{273,273,273,273,0,0,0,2403,0,0,0,0,0,0,0,0,2403,2403,2403,2403,2403,0,0,273,273},
'{273,273,273,273,0,0,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,0,0,273},
'{273,273,273,0,0,0,2403,2403,4005,4005,2403,2403,4005,4005,4005,2403,2403,2403,2403,2403,2403,2403,2403,0,273},
'{273,273,273,0,2403,0,2403,4005,4005,4005,4005,4005,4005,4005,4005,2403,2403,2403,2403,2403,2403,2403,2403,0,273},
'{273,273,0,0,2403,0,2403,4005,4005,4005,4005,4005,4005,4005,4005,4005,2403,2403,2403,0,2403,2403,2403,0,273},
'{273,273,0,2403,2403,0,2403,4005,4005,4005,4005,4005,4005,4005,4005,4005,4005,2403,2403,0,2403,2403,2403,0,273},
'{273,273,0,2403,2403,0,2403,4005,4005,4005,4005,4005,4005,4005,4005,4005,4005,2403,2403,0,2403,2403,2403,0,273},
'{273,273,0,0,2403,0,2403,4005,4005,4005,4005,4005,4005,4005,4005,4005,4005,2403,2403,2403,0,2403,2403,0,273},
'{273,273,273,0,0,0,2403,4005,4005,4005,4005,4005,4005,4005,4005,4005,4005,2403,2403,2403,0,0,0,273,273},
'{273,273,273,273,273,0,0,4005,4005,4005,4005,4005,4005,4005,4005,4005,4005,2403,2403,2403,0,273,273,273,273},
'{273,273,273,273,273,0,0,0,4005,4005,4005,4005,4005,4005,4005,4005,2403,2403,2403,2403,0,273,273,273,273},
'{273,273,273,273,0,2403,2403,0,0,0,4005,4005,4005,4005,2403,2403,2403,2403,2403,2403,0,0,273,273,273},
'{273,273,273,273,0,2403,2403,2403,2403,0,0,0,0,0,2403,2403,2403,2403,2403,2403,2403,0,0,273,273},
'{273,273,273,0,0,2403,2403,2403,2403,2403,2403,0,273,0,2403,2403,2403,2403,2403,2403,2403,2403,0,0,0},
'{273,273,273,0,2403,2403,2403,2403,2403,2403,0,0,273,0,0,2403,2403,2403,2403,2403,2403,2403,0,273,273},
'{273,273,273,0,2403,2403,2403,2403,2403,2403,0,273,273,273,0,0,2403,2403,2403,2403,2403,0,0,273,273},
'{273,273,273,0,0,2403,2403,2403,2403,0,0,273,273,273,273,0,0,2403,2403,2403,0,0,273,273,273},
'{273,273,273,273,0,0,0,0,0,273,273,273,273,273,273,273,0,0,0,0,0,273,273,273,273}
};




parameter bit [11:0] DeadJerryColors1 [29][37] = '{
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,0,0,0,0,273,273,273,273},
'{273,273,273,819,0,0,0,0,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,273,273,273,0,273,273,273,273},
'{273,273,0,0,0,2403,2403,2403,0,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,0,0,273,0,273,273,273,273},
'{273,273,0,0,2403,4005,4005,2403,2403,0,0,273,273,273,273,273,273,0,273,273,273,273,273,273,273,273,273,273,273,273,273,0,0,273,273,273,273},
'{273,0,0,2403,4005,4005,4005,4005,2403,2403,0,273,273,273,273,273,0,0,0,0,0,0,0,0,0,0,273,273,273,0,0,0,273,273,273,273,273},
'{273,0,2403,3989,4005,4005,4005,4005,0,2403,0,0,0,0,0,0,0,2403,2403,2403,2403,2403,2403,2403,2403,0,0,0,0,0,0,0,0,273,273,273,273},
'{273,0,2659,4006,4005,4005,4005,4005,0,2403,2131,2403,2403,2403,2403,2403,0,0,0,0,2403,2403,2403,2659,2659,0,2403,2403,2403,2403,2403,2403,0,0,0,273,273},
'{273,0,2403,4005,4005,4005,4006,0,0,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,0,0,0,2403,2403,2403,0,2403,2403,2403,2403,2403,2403,2403,2403,0,0,273},
'{273,0,2403,4006,4005,4005,0,0,2403,2403,2403,2403,2403,0,0,2403,0,0,2659,2403,2403,0,0,0,0,0,2403,2403,2403,2403,2403,2403,2403,2403,2403,0,273},
'{273,0,2403,2403,0,0,0,2131,2659,2403,2403,2403,2403,0,2403,2403,2403,0,2659,2403,2403,2403,2659,4006,4005,4005,4006,4005,2659,2403,2403,2403,2403,2403,2403,0,273},
'{273,0,2403,2403,2403,2403,2403,2659,2403,2403,2403,2403,0,0,2659,2403,2403,0,0,2403,2659,2659,4005,4005,4005,4005,4005,4005,4005,2403,2403,2403,2403,2403,0,0,273},
'{273,0,0,0,2403,0,0,2659,0,2403,0,2403,0,2403,0,0,2403,2403,0,2403,4005,4005,4005,4005,4005,3618,4005,3618,4005,2659,2403,2403,2403,0,0,273,273},
'{273,273,273,0,0,0,2403,2403,2403,0,2403,2403,0,2403,0,4005,4005,2403,0,2403,4005,4005,4005,4005,3618,3618,3618,4005,4005,4005,0,0,0,0,273,273,273},
'{273,273,273,273,0,2403,2403,2403,0,2403,0,2403,0,2403,0,4005,4005,4005,0,2403,4005,4005,4005,4005,3618,3618,3618,4005,3618,4005,0,0,0,0,273,273,273},
'{273,273,273,273,0,2403,2403,2403,2403,2403,2403,2403,0,4005,0,4005,4005,4005,0,2403,2403,4005,4005,4005,4005,3618,4005,3618,4005,4005,0,0,0,0,0,0,273},
'{273,273,273,273,0,2403,2403,2403,2403,2403,2403,2403,4005,4005,4005,4005,4005,4005,0,2403,2403,4005,4005,4005,4005,4005,3618,4005,4005,3989,0,2403,2403,0,0,0,273},
'{273,273,273,273,0,2403,2403,2403,0,2403,0,2403,4005,4005,0,0,4005,4006,0,2403,4005,4005,4005,4005,4005,4005,4005,4005,3618,0,0,2403,2403,2403,2403,0,273},
'{273,273,273,273,0,2403,2403,2403,2403,0,2403,2403,256,4005,0,3925,4005,0,0,2403,3989,4005,4005,4005,4005,4005,4005,4005,4005,0,2659,2403,2403,2403,2403,0,273},
'{273,273,273,273,0,2659,2403,2659,0,2403,0,2403,0,3733,0,3925,4005,0,2403,2403,2403,3989,3989,3989,3989,3989,4005,4005,0,0,2403,2403,2403,2403,0,0,273},
'{273,273,0,0,0,0,2403,2403,2403,2403,2403,2403,0,3989,0,4005,0,0,0,2403,2403,2403,2403,2403,2403,2403,2403,0,0,2403,2403,2403,0,0,0,273,273},
'{273,0,0,2403,2403,0,0,0,2403,2403,2403,2403,3989,4005,4005,4005,0,273,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,273,273,273,273},
'{273,0,2403,2403,2403,2403,2403,0,0,0,0,0,4005,0,4005,0,0,273,0,0,2403,2403,2403,2403,2931,0,273,273,273,273,273,273,273,273,273,273,273},
'{273,0,0,2403,2403,2403,2403,0,0,273,0,0,0,0,0,0,273,273,273,0,0,2403,2403,2403,2659,0,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,0,0,0,0,0,0,273,273,273,0,273,0,273,273,273,273,273,273,0,0,2403,2403,0,0,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,0,273,0,0,273,273,273,273,273,273,0,0,0,0,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,0,0,273,0,0,273,273,273,273,273,273,0,0,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273}
};




parameter bit [11:0] DeadJerryColors2 [37][29] = '{
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,3822,3822,3822,3822,273,273,273,273,273},
'{273,273,273,273,273,0,0,0,273,273,273,273,273,273,273,273,0,0,0,0,0,0,0,0,273,273,273,273,273},
'{273,273,273,273,0,0,2403,0,0,273,273,273,273,273,273,273,0,2403,2403,2403,2403,2659,2403,0,0,273,273,273,273},
'{273,273,273,273,0,2403,2403,2403,0,273,273,273,273,273,273,0,0,2403,2403,4006,4005,4006,3989,2403,0,0,819,273,273},
'{273,273,273,273,0,2403,2403,2403,0,0,0,0,0,0,0,0,2403,2403,0,4005,4005,4005,4005,4005,2403,0,0,273,273},
'{273,273,273,273,0,2403,2403,0,0,2659,2403,2403,2403,2403,2403,0,0,2403,0,4005,4005,4005,4005,4005,4005,2403,0,273,273},
'{273,273,273,273,0,2403,2403,0,2403,2403,2403,2403,2403,2403,2403,2403,0,2403,0,0,4006,4005,4005,4005,4005,2403,0,273,273},
'{273,273,273,273,0,0,0,0,2403,2659,2403,2403,2403,2403,2403,2403,2403,2659,2131,0,0,4005,4005,4005,2403,2403,0,273,273},
'{273,273,273,273,273,0,0,2403,2403,2403,0,0,2403,2403,2403,0,0,2403,2659,2403,0,0,0,2403,2403,0,0,273,273},
'{273,273,273,273,273,273,0,2403,2403,0,2403,2403,0,2403,0,2403,2403,0,2403,2403,2403,2403,2403,2403,0,0,273,273,273},
'{273,273,273,273,273,0,0,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2131,0,0,0,273,273,273,273},
'{273,273,273,0,0,0,0,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,0,273,273,273,273,273,273},
'{273,0,0,273,273,0,4005,3989,0,0,256,4005,4005,0,0,0,0,0,2403,2403,2403,2403,0,273,273,273,273,273,273},
'{273,273,273,0,0,0,0,4005,3989,3733,4005,4005,4005,4005,2403,2403,2403,0,0,0,2403,2403,0,273,273,273,273,273,273},
'{273,273,0,0,273,0,4005,4005,0,0,0,0,4005,0,0,0,0,2659,2403,0,2403,2403,0,273,273,273,273,273,273},
'{273,273,0,273,273,0,0,4005,4005,4005,4005,0,4005,4005,4005,4005,0,2403,2403,2403,2403,2403,0,273,273,273,273,273,273},
'{273,273,273,273,273,273,0,0,0,4005,4005,4005,4005,4005,4005,4005,2403,2403,2403,0,2403,2659,0,0,0,273,273,273,273},
'{273,273,273,273,273,273,273,273,0,0,0,4006,4005,4005,4005,2403,2403,0,0,0,2403,2659,0,2659,0,273,273,273,273},
'{273,273,273,273,273,273,0,0,0,2403,0,0,0,0,0,0,0,0,2659,2659,2403,2659,0,2659,0,273,273,273,273},
'{273,273,273,273,273,0,0,0,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2403,2659,2659,0,2659,0,273,273,273,273},
'{273,273,273,273,0,0,2403,0,2403,2403,3989,4005,2403,2403,4005,4005,4005,2659,2403,2403,2659,2403,0,2659,0,273,273,273,273},
'{273,273,273,0,0,2403,2403,0,2403,3989,4005,4005,4005,4005,4005,4005,4005,2659,2403,2659,0,0,0,2659,0,273,273,273,273},
'{273,273,0,0,2403,2403,2403,0,2403,3989,4005,4005,4005,4005,4005,4005,4005,4005,2659,2659,0,2403,2403,2659,0,273,273,273,273},
'{273,273,0,0,2403,2403,2403,0,2403,3989,4005,4005,4005,4005,4005,4005,4005,4005,4006,2659,0,2659,2403,2659,0,273,273,273,273},
'{273,273,273,0,0,2659,2931,0,2403,3989,4005,4005,4005,4005,3618,3618,4005,4005,4005,2659,0,2659,2403,2659,0,273,273,273,273},
'{273,273,273,273,0,0,0,0,2403,3989,4005,4005,4005,3618,4005,3618,3618,4005,4005,2659,0,0,0,0,0,273,273,273,273},
'{273,273,273,273,273,273,273,0,2403,4005,4005,4005,4005,4005,3618,4005,4005,4005,4006,2403,2403,2403,0,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,0,0,4005,4005,4005,4005,4005,4005,4005,4005,4005,4005,2403,2403,2403,0,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,0,0,0,4005,4005,4005,4005,4005,4005,4005,4005,2659,2403,2403,2403,0,273,273,0,0,0,273},
'{273,273,273,273,273,273,273,0,2403,0,0,0,3989,4005,4005,4005,2659,2403,2403,2403,2403,2403,0,0,273,0,273,0,273},
'{273,273,273,273,273,273,273,0,2403,2403,2659,0,0,0,0,0,2403,2403,2403,2403,2403,2403,0,0,273,0,273,0,273},
'{273,273,273,273,273,273,273,0,2403,2403,2403,2403,2403,0,273,0,2403,2403,2403,2403,2403,2403,0,0,0,273,273,0,273},
'{273,273,273,273,273,273,273,0,0,2403,2403,2403,2403,0,273,0,2403,2403,2403,2403,2403,0,0,273,0,0,0,0,273},
'{273,273,273,273,273,273,273,273,0,2403,2403,2403,0,0,273,0,0,2403,2403,2403,2403,0,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,0,0,2403,2403,0,273,273,273,0,0,2403,2403,0,0,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,0,0,0,0,273,273,273,273,0,0,0,0,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273}
};






















//Jerry Movement
always_ff @( posedge frame_clk or posedge RESET) begin : Movement_Computation
	begin: Move_Jerry
        if (RESET) begin 
            Jerry_Y_Motion <= 10'd0; //Jerry_Y_Step;
			Jerry_X_Motion <= 10'd0; //Jerry_X_Step;
			Jerry_Y_Pos <= Jerry_Y_Center;
			Jerry_X_Pos <= Jerry_X_Center;
			offscreen <= 0;
        end else begin 
			if(Pause) begin
				Jerry_X_Pos <= Jerry_X_Pos;
				Jerry_Y_Pos <= Jerry_Y_Pos;
			end
			else begin
				//if((Jerry_Y_Pos + Jerry_Y_Motion) <= Jerry_Y_Max + 50 ) begin
					Jerry_Y_Pos <= (Jerry_Y_Pos + Jerry_Y_Motion);  // Update Jerry position
				//end
				if((Jerry_X_Pos + Jerry_X_Motion) <= Jerry_X_Max) begin
					Jerry_X_Pos <= (Jerry_X_Pos + Jerry_X_Motion);
				end

				if(Jerry_Y_Pos > Jerry_Y_Max) // jerry has fallen off of the screen
					offscreen <= 1;
				else
					offscreen <= offscreen;

				
				begin
				if ( (Jerry_Y_Pos + height) > Jerry_Y_Max & (Jerry_Y_Pos + height) < Jerry_Y_Max + 150)  begin// Jerry is at the bottom edge, BOUNCE!
					//Jerry_Y_Pos <= Jerry_Y_Max + height; // disabled so that he can fall off of the screen
					//Jerry_Y_Motion <= (~ (Jerry_Y_Step) + 1'b1);  // 2's complement.
					end
						
				else if ( (Jerry_Y_Pos) > Jerry_Y_Max + 150 )  begin// Jerry is at the top edge, BOUNCE!
					Jerry_Y_Pos <= Jerry_Y_Min;
					//Jerry_Y_Motion <= Jerry_Y_Step;
					end
						
				if ( (Jerry_X_Pos + width) > Jerry_X_Max & (Jerry_X_Pos + width) < Jerry_X_Max + 150)  begin// Jerry is at the Right edge, BOUNCE!
					Jerry_X_Pos <= Jerry_X_Max - width;
					//Jerry_X_Motion <= (~ (Jerry_X_Step) + 1'b1);  // 2's complement.
					end
						
				else if ( (Jerry_X_Pos) > Jerry_X_Max + 150 )  begin// Jerry is at the Left edge, BOUNCE!
					Jerry_X_Pos <= Jerry_X_Min;
					//Jerry_X_Motion <= Jerry_X_Step;
					end
				
				else 
				begin
				//Jerry_Y_Motion <= Jerry_Y_Motion;  // Jerry is somewhere in the middle, don't bounce, just keep moving
				//Jerry_X_Motion <= Jerry_X_Motion;
					
				case (KeyCodes)
					8'd04 : begin
								if(Jerry_X_Pos-width > 0) begin
									Jerry_X_Motion <= -Jerry_X_Step;//A
									Jerry_Y_Motion <= 1;
								end
							end
					8'd80 : begin
								if(Jerry_X_Pos-width > 0) begin
									Jerry_X_Motion <= -Jerry_X_Step;//A
									Jerry_Y_Motion <= 1;
								end
							end
							
					8'd07 : begin
								if(Jerry_X_Pos+(width<<1) < 639) begin
									Jerry_X_Motion <= Jerry_X_Step;//D
									Jerry_Y_Motion <= 1;
								end
							end
					8'd79 : begin
								if(Jerry_X_Pos+(width<<1)  < 639) begin
									Jerry_X_Motion <= Jerry_X_Step;//D
									Jerry_Y_Motion <= 1;
								end
							end

								
					8'd81 : begin
								if(Jerry_Y_Pos+height < 479) begin
									Jerry_Y_Motion <= Jerry_Y_Step + 1;//S
									Jerry_X_Motion <= 0;
								end
							end
					8'd22 : begin
								if(Jerry_Y_Pos+height < 479) begin
									Jerry_Y_Motion <= Jerry_Y_Step + 1;//S
									Jerry_X_Motion <= 0;
								end
							end
								
					8'd26 : begin
								//if(Jerry_Y_Pos-height > 0)begin
									// Jerry_Y_Motion <= (~Jerry_Y_Step + 1);//W
									Jerry_Y_Motion <= 1-Jerry_Y_Step;
									Jerry_X_Motion <= 0;
								//end
							end	  
					8'd82 : begin
								if(Jerry_Y_Pos-height > 0)begin
									Jerry_Y_Motion <= 1-Jerry_Y_Step;//W
									Jerry_X_Motion <= 0;
								end
							end	  
					default: begin 
								Jerry_X_Motion <= 1'b0;
								Jerry_Y_Motion <= 1;
							end
				endcase
				end
				
				end
			end		
		end  
    end
end






endmodule