module entities(
input CLK,
input logic RESET, Pause,
input logic frame_clk,
input logic [1:0] KEY,
input logic [7:0] KeyCodes,
input logic [9:0] DrawX, DrawY, 
input logic [50:0] Game_Counter,
output logic [11:0] ColorE,
output logic Active, Death, inc_score, Boss
);


// local variables


logic [9:0] JerryX, JerryY, JerrywidthEnd, JerryheightEnd;
logic [49:0] KilledJerry; // each bit represents whether the player has been killed by that index of tom
logic [11:0] j0Color, st0Color, st1Color, dt0Color, dt1Color, dt2Color, dt3Color, dt4Color, star0Color, star1Color, oneup0Color, oneup1Color, heart0Color, coin0Color, coin1Color, coin2Color, coin3Color, coin4Color, HZ0Color;
logic j0Active, st0Active, st1Active, dt0Active, dt1Active, dt2Active, dt3Active, dt4Active, star0Active, star1Active, oneup0Active, oneup1Active, heart0Active, coin0Active, coin1Active, coin2Active, coin3Active, coin4Active, HZ0Active;
logic [10:0] StarBoost;
logic switch;
logic [6:0] stindx0, stindy0, stindx1, stindy1,dtindx0, dtindy0, dtindx1, dtindy1, dtindx2, dtindy2, dtindx3, dtindy3, dtindx4, dtindy4, starindx0, starindy0, starindx1, starindy1, oneupindx0, oneupindy0, oneupindx1, oneupindy1, coinindx0, coinindy0, coinindx1, coinindy1, coinindx2, coinindy2, coinindx3, coinindy3, coinindx4, coinindy4;
logic [7:0] HZindx0, HZindy0;
logic [9:0] One_Up;
logic [49:0] CheeseCoin;
logic invincibility;
logic [21:0] TenSeconds;
logic [22:0] FiveSeconds;

assign TenSeconds = Game_Counter[49:28];
assign FiveSeconds = Game_Counter[49:27];



assign switch = Game_Counter[25:24] > 1; // switches every so often
assign invincibility = StarBoost > 0;
assign inc_score = CheeseCoin > 0;



//set priority for entities being drawn here
always_comb begin : Pallete_Priority
	if(j0Active)begin
		ColorE = j0Color;
		Active = j0Active;
	end else if(HZ0Active) begin
		ColorE = HZ0Color;
		Active = HZ0Active;
	end else if(star0Active) begin
		ColorE = star0Color;
		Active = star0Active;
	end else if(star1Active) begin
		ColorE = star1Color;
		Active = star1Active;
	end else if(oneup0Active) begin
		ColorE = oneup0Color;
		Active = oneup0Active;
	end else if(oneup1Active) begin
		ColorE = oneup1Color;
		Active = oneup1Active;
	end else if(coin0Active) begin
		ColorE = coin0Color;
		Active = coin0Active;
	end else if(coin1Active) begin
		ColorE = coin1Color;
		Active = coin1Active;
	end else if(coin2Active) begin
		ColorE = coin2Color;
		Active = coin2Active;
	end else if(coin3Active) begin
		ColorE = coin3Color;
		Active = coin3Active;
	end else if(coin4Active) begin
		ColorE = coin4Color;
		Active = coin4Active;
	end else if(st0Active) begin
		ColorE = st0Color;
		Active = st0Active;
	end else if(st1Active) begin
		ColorE = st1Color;
		Active = st1Active;
	end else if(dt0Active) begin
		ColorE = dt0Color;
		Active = dt0Active;
	end else if(dt1Active) begin
		ColorE = dt1Color;
		Active = dt1Active;
	end else if(dt2Active) begin
		ColorE = dt2Color;
		Active = dt2Active;
	end else if(dt3Active) begin
		ColorE = dt3Color;
		Active = dt3Active;
	end else if(dt4Active) begin
		ColorE = dt4Color;
		Active = dt4Active; 
	end else if(heart0Active) begin
		ColorE = heart0Color;
		Active = heart0Active; 
	end else begin
		ColorE = 0;
		Active = 0;
	end
	
end



Jerry j0(
	.*,
	.active(j0Active),
	.Color(j0Color),
	.offscreen(KilledJerry[0]),
	.dead(Death), // KilledJerry[0]   KilledJerry > 0
	.invincibility(invincibility)
);
//


heart h0(
	.*,
    .heart_active(heart0Active),
    .ColorH(heart0Color),
    .death(Death)
);








Smart_Tom st0(
	.*,
	.spawned(TenSeconds > 3), // 5.37 seconds    TenSeconds > 0
	.Color(st0Color),
	.TomColors1(TomColors1[stindy0][stindx0]),
	.TomColors2(TomColors2[stindy0][stindx0]),
	.indx(stindx0), 
	.indy(stindy0),
	.active(st0Active),
	.JerryActive(j0Active),
	.KilledJerry(KilledJerry[10]), // change after testing
	.Invincible(invincibility),
	.X_Start(20),
	.Y_Start(20),
	.X_Step(2),
	.Y_Step(2)
);

Smart_Tom st1(
	.*,
	.spawned(TenSeconds > 6), // 5.37 seconds    TenSeconds > 0
	.Color(st1Color),
	.TomColors1(TomColors1[stindy1][st1indx1]),
	.TomColors2(TomColors2[stindy1][st1indx1]),
	.indx(stindx1), 
	.indy(stindy1),
	.active(st1Active),
	.JerryActive(j0Active),
	.KilledJerry(KilledJerry[11]), // change after testing
	.Invincible(invincibility),
	.X_Start(380),
	.Y_Start(20),
	.X_Step(2),
	.Y_Step(2)
);



Dumb_Tom dt0(
	.*,
	.spawned(FiveSeconds > 0), // 5.37 seconds    TenSeconds > 0
	.Color(dt0Color),
	.TomColors1(TomColors1[dtindy0][dtindx0]),
	.TomColors2(TomColors2[dtindy0][dtindx0]),
	.indx(dtindx0), 
	.indy(dtindy0),
	.active(dt0Active),
	.JerryActive(j0Active),
	.KilledJerry(KilledJerry[1]),
	.Invincible(invincibility),
	.X_Start(200),
	.Y_Start(20),
	.X_Step(6),
	.Y_Step(3)
);


Dumb_Tom dt1(
	.*,
	.spawned(FiveSeconds > 1), // 5.37 seconds    TenSeconds > 0
	.Color(dt1Color),
	.TomColors1(TomColors1[dtindy1][dtindx1]),
	.TomColors2(TomColors2[dtindy1][dtindx1]),
	.indx(dtindx1), 
	.indy(dtindy1),
	.active(dt1Active),
	.JerryActive(j0Active),
	.KilledJerry(KilledJerry[2]),
	.Invincible(invincibility),
	.X_Start(200),
	.Y_Start(20),
	.X_Step(6),
	.Y_Step(3)
);



Dumb_Tom dt2(
	.*,
	.spawned(TenSeconds > 0), // 5.37 seconds    TenSeconds > 0
	.Color(dt2Color),
	.TomColors1(TomColors1[dtindy2][dtindx2]),
	.TomColors2(TomColors2[dtindy2][dtindx2]),
	.indx(dtindx2), 
	.indy(dtindy2),
	.active(dt2Active),
	.JerryActive(j0Active),
	.KilledJerry(KilledJerry[3]),
	.Invincible(invincibility),
	.X_Start(200),
	.Y_Start(20),
	.X_Step(6),
	.Y_Step(3)
);


Dumb_Tom dt3(
	.*,
	.spawned(TenSeconds > 1), // 5.37 seconds    TenSeconds > 0
	.Color(dt3Color),
	.TomColors1(TomColors1[dtindy3][dtindx3]),
	.TomColors2(TomColors2[dtindy3][dtindx3]),
	.indx(dtindx3), 
	.indy(dtindy3),
	.active(dt3Active),
	.JerryActive(j0Active),
	.KilledJerry(KilledJerry[4]),
	.Invincible(invincibility),
	.X_Start(200),
	.Y_Start(20),
	.X_Step(6),
	.Y_Step(3)
);


Dumb_Tom dt4(
	.*,
	.spawned(TenSeconds > 2), // 5.37 seconds    TenSeconds > 0
	.Color(dt4Color),
	.TomColors1(TomColors1[dtindy4][dtindx4]),
	.TomColors2(TomColors2[dtindy4][dtindx4]),
	.indx(dtindx4), 
	.indy(dtindy4),
	.active(dt4Active),
	.JerryActive(j0Active),
	.KilledJerry(KilledJerry[5]),
	.Invincible(invincibility),
	.X_Start(80),
	.Y_Start(220),
	.X_Step(6),
	.Y_Step(3)
);

Star star0(
	.*,
	.spawned(TenSeconds > 0),
	.Color(star0Color),
	.JerryActive(j0Active),
	.StarColors1(StarColors1[starindy0][starindx0]),
	.StarColors2(StarColors2[starindy0][starindx0]),
	.X_Start(320),
	.Y_Start(5),
	.X_Step(6),
	.Y_Step(3),
	.indx(starindx0), 
	.indy(starindy0),
	.active(star0Active), 
	.StarBoost(StarBoost[0])
);
One_UP up0(
	.*,
	.spawned(TenSeconds > 1),
	.JerryActive(j0Active),
	.One_UPColors1(OneUpColors1[oneupindy0][oneupindx0]),
	.One_UPColors2(OneUpColors2[oneupindy0][oneupindx0]), 
	.X_Start(320),
	.Y_Start(5),
	.X_Step(1),
	.Y_Step(1),
	.Color(oneup0Color),
	.indx(oneupindx0), 
	.indy(oneupindy0),
	.active(oneup0Active), 
	.One_Up(One_Up[0])
);

Star star1(
	.*,
	.spawned(TenSeconds > 3),
	.Color(star1Color),
	.JerryActive(j0Active),
	.StarColors1(StarColors1[starindy1][starindx1]),
	.StarColors2(StarColors2[starindy1][starindx1]),
	.X_Start(320),
	.Y_Start(5),
	.X_Step(6),
	.Y_Step(3),
	.indx(starindx1), 
	.indy(starindy1),
	.active(star1Active), 
	.StarBoost(StarBoost[1])
);
One_UP up1(
	.*,
	.spawned(TenSeconds > 4),
	.JerryActive(j0Active),
	.One_UPColors1(OneUpColors1[oneupindy1][oneupindx1]),
	.One_UPColors2(OneUpColors2[oneupindy1][oneupindx1]), 
	.X_Start(320),
	.Y_Start(5),
	.X_Step(2),
	.Y_Step(2),
	.Color(oneup1Color),
	.indx(oneupindx1), 
	.indy(oneupindy1),
	.active(oneup1Active), 
	.One_Up(One_Up[1])
);






CheeseCoin coin0(
	.*,
	.spawned(FiveSeconds > 1),
	.JerryActive(j0Active),
	.CheeseCoinColors1(CheeseCoinColors1[coinindy0][coinindx0]),
	.CheeseCoinColors2(CheeseCoinColors2[coinindy0][coinindx0]), 
	.X_Start(320),
	.Y_Start(5),
	.X_Step(0),
	.Y_Step(Game_Counter[39:30]),
	.Color(coin0Color),
	.indx(coinindx0), 
	.indy(coinindy0),
	.active(coin0Active), 
	.CheeseCoin(CheeseCoin[0])
);


CheeseCoin coin1(
	.*,
	.spawned(FiveSeconds > 2),
	.JerryActive(j0Active),
	.CheeseCoinColors1(CheeseCoinColors1[coinindy1][coinindx1]),
	.CheeseCoinColors2(CheeseCoinColors2[coinindy1][coinindx1]), 
	.X_Start(30),
	.Y_Start(5),
	.X_Step(0),
	.Y_Step(Game_Counter[39:30]),
	.Color(coin1Color),
	.indx(coinindx1), 
	.indy(coinindy1),
	.active(coin1Active), 
	.CheeseCoin(CheeseCoin[1])
);


CheeseCoin coin2(
	.*,
	.spawned(FiveSeconds > 3),
	.JerryActive(j0Active),
	.CheeseCoinColors1(CheeseCoinColors1[coinindy2][coinindx2]),
	.CheeseCoinColors2(CheeseCoinColors2[coinindy2][coinindx2]), 
	.X_Start(180),
	.Y_Start(5),
	.X_Step(0),
	.Y_Step(Game_Counter[39:30]),
	.Color(coin2Color),
	.indx(coinindx2), 
	.indy(coinindy2),
	.active(coin2Active), 
	.CheeseCoin(CheeseCoin[2])
);


CheeseCoin coin3(
	.*,
	.spawned(FiveSeconds > 4),
	.JerryActive(j0Active),
	.CheeseCoinColors1(CheeseCoinColors1[coinindy3][coinindx3]),
	.CheeseCoinColors2(CheeseCoinColors2[coinindy3][coinindx3]), 
	.X_Start(460),
	.Y_Start(5),
	.X_Step(0),
	.Y_Step(Game_Counter[39:30]),
	.Color(coin3Color),
	.indx(coinindx3), 
	.indy(coinindy3),
	.active(coin3Active), 
	.CheeseCoin(CheeseCoin[3])
);


CheeseCoin coin4(
	.*,
	.spawned(FiveSeconds > 5),
	.JerryActive(j0Active),
	.CheeseCoinColors1(CheeseCoinColors1[coinindy4][coinindx4]),
	.CheeseCoinColors2(CheeseCoinColors2[coinindy4][coinindx4]), 
	.X_Start(580),
	.Y_Start(5),
	.X_Step(0),
	.Y_Step(Game_Counter[39:30]),
	.Color(coin4Color),
	.indx(coinindx4), 
	.indy(coinindy4),
	.active(coin4Active), 
	.CheeseCoin(CheeseCoin[4])
);





























always_ff @( posedge CLK or posedge RESET ) begin : BossButton
	if(RESET)
		Boss <= 0;
	else begin
		if(KEY[1])
			Boss <= Boss;
		else
			Boss <= 1;
	end
end



HZ hz0( // the boss himself
	.*,
	.spawned(Boss), // 5.37 seconds    
	.Color(HZ0Color),
	.HZColors1(HZColors1[HZindy0][HZindx0]),
	.HZColors2(HZColors2[HZindy0][HZindx0]),
	.indx(HZindx0), 
	.indy(HZindy0),
	.active(HZ0Active),
	.Invincible(invincibility),
	.JerryActive(j0Active),
	.KilledJerry(KilledJerry[49]), // change after testing
	.X_Start(20),
	.Y_Start(20),
	.X_Step(2),
	.Y_Step(2)
);





//Tom definition
parameter bit [11:0] TomColors1 [40][40] = '{
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,0,0,0,0,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,4095,4095,4095,0,0,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,0,0,0,273,273,273,273,273,0,0,4095,4095,4095,2201,0,0,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,0,0,0,273,273,273,273,273,0,0,0,4026,0,273,273,273,273,273,273,273,0,0,0,0,2201,2201,0,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,0,0,0,273,273,273,0,0,2201,0,4026,0,273,273,273,273,273,273,273,273,273,273,0,0,2201,2201,0,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,0,0,0,0,0,0,0,2201,0,4026,4026,0,273,273,273,273,273,273,273,273,273,273,273,0,0,2201,0,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,0,2201,2201,2201,2201,2201,2201,2201,0,4026,0,273,273,273,273,273,273,273,273,273,273,273,273,273,0,2201,0,273,273,273},
'{273,273,273,273,273,273,273,273,273,0,0,0,2201,2201,2201,2201,0,0,2201,2201,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2201,0,273,273,273},
'{273,273,273,273,273,273,273,273,0,0,2201,0,0,2201,2201,0,0,2201,2201,2201,0,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,0,273,273,273},
'{273,273,273,273,273,273,273,273,0,2201,2201,4073,0,2201,2201,0,4073,2201,2201,2201,0,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,0,273,273,273},
'{273,273,273,273,273,273,0,0,0,2201,2201,4095,4095,4095,4095,4095,2201,2201,2201,0,0,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,0,273,273,273},
'{273,273,273,0,0,0,0,2201,0,2201,4095,4095,0,0,4095,4095,4095,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,0,0,273,273},
'{273,273,273,0,4095,2201,2201,2201,2201,0,0,4095,4095,4095,4095,4095,4095,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,0,273,273},
'{273,273,0,0,4095,4095,0,0,0,0,0,0,4095,4095,4095,4095,0,0,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,0,273,273},
'{273,273,0,4095,4095,0,0,273,273,273,273,0,0,0,0,0,0,2201,2201,2201,2201,4095,4095,4095,4095,4095,4095,4095,4095,2201,2201,2201,2201,2201,2201,2201,2201,0,0,273},
'{273,273,0,0,0,0,273,273,273,273,273,273,273,0,0,0,2201,2201,2201,2201,0,0,0,0,0,0,0,0,4095,4095,2201,2201,2201,2201,2201,2201,2201,2201,0,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,0,0,2201,2201,2201,2201,2201,0,0,273,273,273,273,0,0,0,0,4095,2201,2201,2201,2201,2201,2201,2201,2201,0,273},
'{273,273,273,273,273,273,273,273,273,273,0,0,0,2201,2201,2201,2201,0,0,0,273,273,273,273,273,0,2201,2201,0,0,0,0,2201,2201,2201,2201,2201,2201,0,273},
'{273,273,273,273,273,273,273,273,0,0,0,4095,2201,2201,2201,2201,0,0,273,273,273,273,273,273,0,0,2201,2201,2201,2201,0,0,0,2201,2201,2201,2201,0,0,273},
'{273,273,273,273,273,273,273,273,0,4095,4095,4095,4095,4095,2201,0,0,273,273,273,273,273,273,0,0,2201,2201,2201,2201,2201,0,273,0,0,2201,2201,2201,0,273,273},
'{273,273,273,273,273,273,273,273,0,4095,4095,4095,4095,0,0,0,273,273,273,273,273,0,0,0,2201,2201,2201,2201,0,0,0,0,0,2201,2201,2201,2201,0,273,273},
'{273,273,273,273,273,273,273,273,273,0,0,0,0,0,273,273,273,273,273,0,0,0,4095,4095,2201,2201,0,0,0,4095,4095,4095,2201,2201,2201,0,0,0,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,4095,4095,4095,4095,4095,0,0,0,4095,4095,4095,4095,4095,2201,0,0,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,0,0,0,0,0,0,273,0,0,0,0,0,0,0,0,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273}
};


parameter bit [11:0] TomColors2 [40][40] = '{
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,0,0,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,0,4095,0,0,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,4095,4095,0,0,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,4095,4095,4095,0,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,0,0,0,273,273,273,273,273,273,273,273,273,0,0,4095,4095,0,273,273,273},
'{273,273,273,273,273,273,273,273,273,0,0,0,273,273,273,273,273,0,0,0,4026,0,273,273,273,273,273,273,273,273,273,273,273,0,2201,2201,0,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,0,0,0,273,273,273,0,0,2201,0,4026,0,273,273,273,273,273,273,273,273,273,273,273,0,0,2201,0,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,0,0,0,0,0,0,0,2201,0,4026,4026,0,273,273,273,273,273,273,273,273,273,273,273,273,0,2201,0,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,0,2201,2201,2201,2201,2201,2201,2201,0,4026,0,273,273,273,273,273,273,273,273,273,273,273,273,273,0,2201,0,273,273,273},
'{273,273,273,273,273,273,273,273,273,0,0,0,2201,2201,2201,2201,0,0,2201,2201,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2201,0,273,273,273},
'{273,273,273,273,273,273,273,273,0,0,2201,0,0,2201,2201,0,0,2201,2201,2201,0,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,0,273,273,273},
'{273,273,0,0,0,0,0,0,0,2201,2201,4073,0,2201,2201,0,4073,2201,2201,2201,0,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,0,273,273,273},
'{273,0,0,4095,4095,4095,2201,2201,0,2201,2201,4095,4095,4095,4095,4095,2201,2201,2201,0,0,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,0,273,273,273},
'{273,0,0,0,0,0,2201,2201,0,2201,4095,4095,0,0,4095,4095,4095,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,0,0,273,273},
'{273,273,273,273,273,0,0,0,0,0,0,4095,4095,4095,4095,4095,4095,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,0,273,273},
'{273,273,273,273,273,273,273,273,273,273,0,0,4095,4095,4095,4095,0,0,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,2201,0,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,0,0,0,0,0,0,2201,2201,2201,2201,4095,4095,4095,4095,4095,4095,4095,4095,2201,2201,2201,2201,2201,2201,2201,2201,0,0,273},
'{273,273,273,273,273,273,273,273,273,0,0,0,0,2201,2201,2201,2201,2201,2201,0,0,0,0,0,0,0,0,0,0,0,2201,2201,2201,2201,2201,2201,2201,2201,0,273},
'{273,273,273,273,273,273,0,0,0,0,4095,2201,2201,2201,2201,2201,2201,2201,0,0,273,273,273,273,273,0,0,2201,2201,0,0,0,2201,2201,2201,2201,2201,2201,0,273},
'{273,273,273,273,273,273,0,4095,4095,4095,4095,4095,2201,2201,2201,2201,0,0,0,273,273,273,273,0,273,0,2201,2201,2201,2201,2201,0,2201,2201,2201,2201,2201,2201,0,273},
'{273,273,273,273,273,273,0,0,4095,4095,4095,4095,2201,2201,2201,0,0,273,273,273,273,273,273,273,273,0,2201,2201,2201,2201,0,0,0,2201,2201,2201,2201,2201,0,273},
'{273,273,273,273,273,273,273,0,0,0,0,0,0,0,0,0,273,273,273,273,273,273,273,273,273,273,2201,2201,2201,2201,0,273,0,2201,2201,2201,2201,2201,0,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,2201,2201,2201,2201,0,273,273,0,2201,2201,2201,2201,2201,0,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,2201,2201,2201,2201,0,273,273,0,2201,2201,2201,2201,2201,0,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,2201,2201,2201,0,0,273,273,0,0,2201,2201,2201,2201,0,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,0,0,4095,2201,2201,0,273,273,273,273,0,0,2201,2201,2201,0,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,0,4095,4095,4095,4095,0,0,273,273,273,273,273,0,4095,4095,4095,0,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,0,4095,4095,4095,4095,0,0,273,273,273,273,273,0,0,4095,4095,0,0,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,0,0,0,0,0,273,273,273,273,273,273,0,4095,4095,4095,0,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,0,0,0,0,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273}
};






parameter bit [11:0] StarColors1 [35][35] = '{
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,3696,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,3696,3696,3696,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,3696,4064,3696,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,3696,4064,4064,4064,3696,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,3696,4064,4064,4064,3696,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,3696,4064,4064,4064,4064,4064,3696,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,3696,4064,4064,4064,4064,4064,3696,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,3696,4064,4064,4064,4064,4064,4064,4064,3696,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,3696,4064,4064,4064,4064,4064,4064,4064,3696,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,4064,4064,4064,4048,4064,4048,4064,4064,4064,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,273,273},
'{273,273,3696,3696,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,3696,3696,273,273},
'{273,273,273,3696,3696,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,3696,3696,273,273,273},
'{273,273,273,273,3696,3696,4064,4064,4064,4064,4064,4064,4064,4064,3696,3696,4064,4064,4064,3696,3696,4064,4064,4064,4064,4064,4064,4064,4064,3696,3696,273,273,273,273},
'{273,273,273,273,273,3696,3696,4064,4064,4064,4064,4064,4064,4064,3696,3696,4064,4064,4064,3696,3696,4064,4064,4064,4064,4064,4064,4064,3696,3696,273,273,273,273,273},
'{273,273,273,273,273,273,3696,3696,4064,4064,4064,4064,4064,4064,3696,3696,4064,4064,4064,3696,3696,4064,4064,4064,4064,4064,4064,3696,3696,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,3696,3696,4064,4064,4064,4064,4064,3696,3696,4064,4064,4064,3696,3696,4064,4064,4064,4064,4064,3696,3696,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,3696,3696,4064,4064,4064,4064,3696,3696,4064,4064,4064,3696,3696,4064,4064,4064,4064,3696,3696,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,3696,3696,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,3696,3696,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,3696,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,3696,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,3696,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,3696,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,3696,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,3696,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,3696,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,3696,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,3696,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,3696,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,3696,4064,4064,4064,4064,4064,4064,4064,4064,3696,3696,3696,4064,4064,4064,4064,4064,4064,4064,4064,3696,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,3696,4064,4064,4064,4064,4064,4064,4064,4064,3696,3696,273,3696,3696,4064,4064,4064,4064,4064,4064,4064,4064,3696,273,273,273,273,273,273},
'{273,273,273,273,273,273,3696,4064,4064,4064,4064,4064,4064,3696,3696,3696,273,273,273,3696,3696,3696,4064,4064,4064,4064,4064,4064,3696,273,273,273,273,273,273},
'{273,273,273,273,273,3696,4064,4064,4064,4064,4064,3696,3696,3696,273,273,273,273,273,273,273,3696,3696,3696,4064,4064,4064,4064,4064,3696,273,273,273,273,273},
'{273,273,273,273,3696,4064,4064,4064,4064,3696,3696,3696,273,273,273,273,273,273,273,273,273,273,273,3696,3696,3696,4064,4064,4064,4064,3696,273,273,273,273},
'{273,273,273,273,3696,4064,4064,3696,3696,3696,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,3696,3696,3696,4064,4064,3696,273,273,273,273},
'{273,273,273,3696,4064,3696,3696,3696,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,3696,3696,3696,4064,3696,273,273,273},
'{273,273,273,3696,3696,3696,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,3696,3696,3696,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273}
};







parameter bit [11:0] StarColors2 [35][35] = '{
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,4064,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,4064,4064,4064,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,4064,3696,4064,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,4064,3696,3696,3696,4064,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,4064,3696,3696,3696,4064,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,4064,3696,3696,3696,3696,3696,4064,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,4064,3696,3696,3696,3696,3696,4064,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,4064,3696,3696,3696,3696,3696,3696,3696,4064,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,4064,3696,3696,3696,3696,3696,3696,3696,4064,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,3424,3696,3696,3696,3696,3696,3696,3696,3424,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,273,273},
'{273,273,4064,4064,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,4064,4064,273,273},
'{273,273,273,4064,4064,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,4064,4064,273,273,273},
'{273,273,273,273,4064,4064,3696,3696,3696,3696,3696,3696,3696,3696,4064,4064,3696,3696,3696,4064,4064,3696,3696,3696,3696,3696,3696,3696,3696,4064,4064,273,273,273,273},
'{273,273,273,273,273,4064,4064,3696,3696,3696,3696,3696,3696,3696,4064,4064,3696,3696,3696,4064,4064,3696,3696,3696,3696,3696,3696,3696,4064,4064,273,273,273,273,273},
'{273,273,273,273,273,273,4064,4064,3696,3696,3696,3696,3696,3696,4064,4064,3696,3696,3696,4064,4064,3696,3696,3696,3696,3696,3696,4064,4064,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,4064,4064,3696,3696,3696,3696,3696,4064,4064,3696,3696,3696,4064,4064,3696,3696,3696,3696,3696,4064,4064,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,4064,4064,3696,3696,3696,3696,4064,4064,3696,3696,3696,4064,4064,3696,3696,3696,3696,4064,4064,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,4064,4064,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,4064,4064,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,4064,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,4064,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,4064,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,4064,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,4064,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,4064,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,4064,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,4064,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,4064,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,3696,4064,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,4064,3696,3696,3696,3696,3696,3696,3696,3696,4064,4064,4064,3696,3696,3696,3696,3696,3696,3696,3696,4064,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,4064,3696,3696,3696,3696,3696,3696,3696,3696,4064,4064,273,4064,4064,3696,3696,3696,3696,3696,3696,3696,3696,4064,273,273,273,273,273,273},
'{273,273,273,273,273,273,4064,3696,3696,3696,3696,3696,3696,4064,4064,4064,273,273,273,4064,4064,4064,3696,3696,3696,3696,3696,3696,4064,273,273,273,273,273,273},
'{273,273,273,273,273,4064,3696,3696,3696,3696,3696,4064,4064,4064,273,273,273,273,273,273,273,4064,4064,4064,3696,3696,3696,3696,3696,4064,273,273,273,273,273},
'{273,273,273,273,4064,3696,3696,3696,3696,4064,4064,4064,273,273,273,273,273,273,273,273,273,273,273,4064,4064,4064,3696,3696,3696,3696,4064,273,273,273,273},
'{273,273,273,273,4064,3696,3696,4064,4064,4064,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,4064,4064,4064,3696,3696,4064,273,273,273,273},
'{273,273,273,4064,3696,4064,4064,4064,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,4064,4064,4064,3696,4064,273,273,273},
'{273,273,273,4064,4064,4064,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,4064,4064,4064,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273}
};





parameter bit [11:0] OneUpColors1 [25][25] = '{
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,0,0,0,0,0,0,0,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,0,0,0,4095,146,146,146,4095,0,0,0,273,273,273,273,273,273,273},
'{273,273,273,273,273,0,0,0,4095,4095,4095,146,146,146,4095,4095,4095,0,0,0,273,273,273,273,273},
'{273,273,273,273,0,0,4095,4095,4095,4095,4095,146,146,146,4095,4095,4095,4095,4095,0,0,273,273,273,273},
'{273,273,273,0,0,146,4095,4095,4095,4095,146,146,146,146,146,146,4095,4095,4095,146,0,0,273,273,273},
'{273,273,273,0,4095,146,146,146,4095,4095,4095,4095,4095,4095,4095,146,146,146,146,146,4095,0,273,273,273},
'{273,273,0,0,4095,4095,146,146,4095,4095,4095,4095,4095,4095,4095,4095,4095,146,146,4095,4095,0,0,273,273},
'{273,273,0,4095,4095,4095,146,146,4095,4095,4095,4095,4095,4095,4095,4095,4095,146,146,4095,4095,4095,0,273,273},
'{273,273,0,4095,4095,4095,146,146,4095,4095,4095,4095,4095,4095,4095,4095,4095,146,146,4095,4095,4095,0,273,273},
'{273,273,0,4095,4095,4095,146,146,4095,4095,4095,4095,4095,4095,4095,4095,4095,146,146,4095,4095,4095,0,273,273},
'{273,273,0,4095,4095,146,146,146,4095,4095,4095,4095,4095,4095,4095,4095,4095,146,146,146,4095,4095,0,273,273},
'{273,273,0,146,146,146,146,146,146,146,4095,4095,4095,4095,4095,146,146,146,146,146,146,146,0,273,273},
'{273,273,0,146,146,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,146,146,0,273,273},
'{273,0,0,0,0,0,4095,4095,4095,0,0,4095,4095,4095,0,0,4095,4095,4095,0,0,0,0,0,273},
'{273,273,273,0,0,4095,4095,4095,4095,0,0,4095,4095,4095,0,0,4095,4095,4095,4095,0,0,273,273,273},
'{273,273,273,273,0,4095,4095,4095,4095,0,0,4095,4095,4095,0,0,4095,4095,4095,4095,0,273,273,273,273},
'{273,273,273,273,0,0,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,0,0,273,273,273,273},
'{273,273,273,273,273,0,0,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,0,0,273,273,273,273,273},
'{273,273,273,273,273,273,0,0,0,0,0,0,0,0,0,0,0,0,0,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273}
};




parameter bit [11:0] OneUpColors2 [25][25] = '{
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,0,0,0,0,0,0,0,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,0,0,0,4095,146,146,146,4095,0,0,0,273,273,273,273,273,273,273},
'{273,273,273,273,273,0,0,0,4095,4095,4095,146,146,146,4095,4095,4095,0,0,0,273,273,273,273,273},
'{273,273,273,273,0,0,4095,4095,4095,4095,4095,146,146,146,4095,4095,4095,4095,4095,0,0,273,273,273,273},
'{273,273,273,0,0,146,4095,4095,4095,146,146,146,146,146,146,146,4095,4095,4095,146,0,0,273,273,273},
'{273,273,273,0,4095,146,146,146,146,146,4095,4095,4095,4095,4095,146,146,146,146,146,4095,0,273,273,273},
'{273,273,0,0,4095,4095,146,146,4095,4095,4095,4095,4095,4095,4095,4095,4095,146,146,4095,4095,0,0,273,273},
'{273,273,0,4095,4095,4095,146,146,4095,4095,4095,4095,4095,4095,4095,4095,4095,146,146,4095,4095,4095,0,273,273},
'{273,273,0,4095,4095,4095,146,146,4095,4095,4095,4095,4095,4095,4095,4095,4095,146,146,4095,4095,4095,0,273,273},
'{273,0,0,4095,4095,4095,146,146,4095,4095,4095,4095,4095,4095,4095,4095,4095,146,146,4095,4095,4095,0,273,273},
'{273,0,0,4095,4095,146,146,146,4095,4095,4095,4095,4095,4095,4095,4095,4095,146,146,146,4095,4095,0,273,273},
'{273,273,0,146,146,146,146,146,146,146,4095,4095,4095,4095,4095,146,146,146,146,146,146,146,0,273,273},
'{273,273,0,146,146,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,146,146,0,273,273},
'{273,0,0,0,0,0,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,0,0,0,0,273,273},
'{273,273,273,0,0,4095,4095,4095,0,0,0,4095,4095,4095,0,0,0,4095,4095,4095,0,0,273,273,273},
'{273,273,273,273,0,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,0,273,273,273,273},
'{273,273,273,273,0,0,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,0,0,273,273,273,273},
'{273,273,273,273,273,0,0,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,4095,0,0,273,273,273,273,273},
'{273,273,273,273,273,273,0,0,0,0,0,0,0,0,0,0,0,0,0,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273}
};





parameter bit [11:0] CheeseCoinColors1 [25][32] = '{
'{273,273,273,273,273,273,273,273,273,0,0,0,0,0,0,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,0,4064,4064,4064,4064,4064,4064,0,0,0,0,0,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,0,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,0,0,0,0,0,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,0,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,0,0,0,273,273,273,273},
'{273,273,273,273,273,273,0,4064,4064,4064,4064,4064,0,0,0,4064,4064,4064,4064,4064,4064,0,0,0,0,4064,4064,0,0,273,273,273},
'{273,273,273,273,273,0,4064,4064,4064,4064,4064,0,4023,4023,4023,0,4064,4064,0,0,0,4064,4064,4064,4064,4064,4064,4064,0,273,273,273},
'{273,273,273,273,0,4064,4064,4064,4064,4064,0,4023,4023,4023,4023,4023,0,0,0,4064,4064,4064,4064,4064,4064,4064,0,0,0,273,273,273},
'{273,273,273,0,4064,4064,4064,0,0,0,0,4023,4023,4023,4023,4023,0,4064,4064,4064,4064,4064,4064,4064,4064,0,4023,0,273,273,273,273},
'{273,273,0,4064,0,0,0,4064,4064,4064,0,4023,4023,4023,4023,4023,0,4064,4064,0,4064,4064,4064,4064,4064,0,4023,0,273,273,273,273},
'{273,273,0,0,4064,4064,4064,4064,4064,4064,4064,0,4023,4023,4023,0,4064,4064,0,4023,0,4064,4064,4064,4064,4064,0,0,0,273,273,273},
'{273,0,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,0,0,0,4064,4064,4064,4064,0,4064,4064,4064,4064,4064,4064,4064,4064,0,273,273,273},
'{273,0,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,0,0,4064,4064,4064,4064,4064,4064,4064,4064,0,0,0,273,273,273},
'{273,0,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,0,4023,4023,0,4064,4064,4064,4064,4064,4064,0,4023,4023,0,273,273,273},
'{273,0,0,0,0,4064,4064,4064,4064,0,4064,4064,4064,4064,4064,4064,0,0,4064,4064,4064,4064,4064,4064,0,4023,4023,0,273,273,273,273},
'{273,273,0,4023,0,4064,4064,4064,0,4023,0,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,0,4023,4023,0,273,273,273,273},
'{273,273,0,4023,4023,0,4064,4064,4064,0,4064,4064,4064,4064,0,0,0,4064,4064,4064,4064,4064,4064,4064,0,4023,4023,0,0,273,273,273},
'{273,273,273,0,4023,0,4064,4064,4064,4064,4064,4064,4064,0,4023,4023,4023,0,4064,4064,4064,4064,4064,4064,4064,0,4023,4023,0,273,273,273},
'{273,273,0,4023,4023,0,4064,4064,4064,4064,4064,4064,0,4023,4023,4023,4023,4023,0,4064,4064,4064,4064,4064,4064,4064,0,0,0,273,273,273},
'{273,273,0,4023,0,4064,4064,4064,4064,4064,4064,0,4023,4023,4023,4023,4023,4023,4023,0,4064,4064,4064,4064,0,0,0,0,273,273,273,273},
'{273,0,0,0,0,4064,4064,4064,4064,4064,4064,0,4023,4023,0,0,0,4023,0,4023,0,0,0,0,273,273,273,273,273,273,273,273},
'{273,0,4064,4064,4064,4064,4064,4064,4064,4064,4064,0,4023,0,273,273,273,0,0,0,0,273,273,273,273,273,273,273,273,273,273,273},
'{273,0,4064,4064,4064,4064,4064,4064,4064,4064,4064,4064,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,0,4064,4064,4064,4064,4064,4064,0,0,0,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,0,0,0,0,0,0,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273}
};





parameter bit [11:0] CheeseCoinColors2 [25][32] = '{
'{273,273,273,273,273,273,273,273,273,0,0,0,0,0,0,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,0,4023,4023,4023,4023,4023,4023,0,0,0,0,0,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,0,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,0,0,0,0,0,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,0,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,0,0,0,273,273,273,273},
'{273,273,273,273,273,273,0,4023,4023,4023,4023,4023,0,0,0,4023,4023,4023,4023,4023,4023,0,0,0,0,4023,4023,0,0,273,273,273},
'{273,273,273,273,273,0,4023,4023,4023,4023,4023,0,4064,4064,4064,0,4023,4023,0,0,0,4023,4023,4023,4023,4023,4023,4023,0,273,273,273},
'{273,273,273,273,0,4023,4023,4023,4023,4023,0,4064,4064,4064,4064,4064,0,0,0,4023,4023,4023,4023,4023,4023,4023,0,0,0,273,273,273},
'{273,273,273,0,4023,4023,4023,0,0,0,0,4064,4064,4064,4064,4064,0,4023,4023,4023,4023,4023,4023,4023,4023,0,4064,0,273,273,273,273},
'{273,273,0,4023,0,0,0,4023,4023,4023,0,4064,4064,4064,4064,4064,0,4023,4023,0,4023,4023,4023,4023,4023,0,4064,0,273,273,273,273},
'{273,273,0,0,4023,4023,4023,4023,4023,4023,4023,0,4064,4064,4064,0,4023,4023,0,4064,0,4023,4023,4023,4023,4023,0,0,0,273,273,273},
'{273,0,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,0,0,0,4023,4023,4023,4023,0,4023,4023,4023,4023,4023,4023,4023,4023,0,273,273,273},
'{273,0,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,0,0,4023,4023,4023,4023,4023,4023,4023,4023,0,0,0,273,273,273},
'{273,0,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,0,4064,4064,0,4023,4023,4023,4023,4023,4023,0,4064,4064,0,273,273,273},
'{273,0,0,0,0,4023,4023,4023,4023,0,4023,4023,4023,4023,4023,4023,0,0,4023,4023,4023,4023,4023,4023,0,4064,4064,0,273,273,273,273},
'{273,273,0,4064,0,4023,4023,4023,0,4064,0,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,0,4064,4064,0,273,273,273,273},
'{273,273,0,4064,4064,0,4023,4023,4023,0,4023,4023,4023,4023,0,0,0,4023,4023,4023,4023,4023,4023,4023,0,4064,4064,0,0,273,273,273},
'{273,273,273,0,4064,0,4023,4023,4023,4023,4023,4023,4023,0,4064,4064,4064,0,4023,4023,4023,4023,4023,4023,4023,0,4064,4064,0,273,273,273},
'{273,273,0,4064,4064,0,4023,4023,4023,4023,4023,4023,0,4064,4064,4064,4064,4064,0,4023,4023,4023,4023,4023,4023,4023,0,0,0,273,273,273},
'{273,273,0,4064,0,4023,4023,4023,4023,4023,4023,0,4064,4064,4064,4064,4064,4064,4064,0,4023,4023,4023,4023,0,0,0,0,273,273,273,273},
'{273,0,0,0,0,4023,4023,4023,4023,4023,4023,0,4064,4064,0,0,0,4064,0,4064,0,0,0,0,273,273,273,273,273,273,273,273},
'{273,0,4023,4023,4023,4023,4023,4023,4023,4023,4023,0,4064,0,273,273,273,0,0,0,0,273,273,273,273,273,273,273,273,273,273,273},
'{273,0,4023,4023,4023,4023,4023,4023,4023,4023,4023,4023,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,0,4023,4023,4023,4023,4023,4023,0,0,0,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,0,0,0,0,0,0,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273}
};









parameter bit [11:0] HZColors1 [170][125] = '{
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,4095,2457,2457,2457,2457,2458,2458,2458,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2191,2459,2458,2185,2457,2457,2457,2185,2185,2184,1912,1912,2184,2184,2184,2185,2458,4095,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,2184,2184,2184,2185,2185,2185,2184,1912,1912,1912,1912,1912,1911,1639,1638,1638,1639,1639,1639,1911,2184,2185,2458,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2730,2457,2185,2184,1912,1639,1639,1639,1639,1911,1911,1639,1638,1638,1639,1638,1638,1366,1365,1093,1093,1365,1365,1365,1366,1639,1912,2185,2457,2458,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2186,2457,2185,2185,2184,1912,1911,1638,1366,1366,1366,1366,1366,1366,1366,1365,1365,1365,1365,1093,1093,1092,820,820,820,1092,1092,1093,1366,1639,1911,2184,2185,2185,2185,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2457,2185,2185,2185,2184,1912,1911,1911,1639,1638,1365,1093,1092,1092,1092,1092,1093,1092,820,820,820,820,820,820,819,547,547,547,547,547,819,1092,1365,1638,1911,1911,1912,1912,2185,2457,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2457,2185,2184,1912,1911,1639,1639,1638,1638,1366,1365,1365,1092,820,819,819,819,819,820,819,547,547,547,547,547,547,546,546,274,274,274,546,547,819,1092,1365,1638,1638,1638,1639,1912,2184,2457,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,2185,2184,1912,1911,1639,1638,1366,1365,1093,1093,1093,1092,1092,1092,819,547,547,546,546,547,547,546,546,546,546,546,546,546,530,274,274,274,274,274,546,547,819,1092,1365,1365,1365,1365,1638,1911,1912,2185,2457,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,2185,2184,1911,1639,1638,1366,1365,1093,820,820,819,819,819,819,819,819,547,546,530,274,274,274,530,274,274,274,274,274,274,274,274,274,274,274,274,274,274,546,547,819,1092,1092,820,1092,1093,1366,1639,1912,2184,2185,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1912,1911,1638,1366,1365,1093,1093,1092,820,819,547,546,546,546,546,546,546,546,274,274,274,274,274,274,274,274,274,274,274,274,274,274,274,274,274,274,274,274,274,546,547,819,819,819,819,820,1092,1365,1638,1639,1911,1912,2184,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1911,1638,1365,1093,1092,820,819,819,819,547,546,274,274,274,274,274,274,274,274,274,274,274,274,274,274,257,1,1,1,1,274,274,274,274,274,1,1,257,274,274,274,546,546,546,546,546,547,819,820,1093,1365,1365,1638,1911,1912,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1911,1638,1365,1092,820,819,547,547,547,546,546,274,274,274,274,274,274,274,274,274,274,274,274,274,274,257,1,1,1,1,1,274,274,274,274,257,1,1,1,274,274,274,274,274,274,274,274,530,546,547,820,820,1092,1093,1366,1638,1912,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1912,1638,1365,1092,819,547,546,546,274,274,530,274,274,274,274,274,274,274,274,274,274,274,274,274,274,1,1,1,257,1,1,1,257,274,274,274,1,1,1,1,1,274,274,274,274,274,274,274,274,274,546,546,547,547,819,1092,1365,1638,1912,2187,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1912,1638,1365,1092,819,547,546,274,274,274,274,274,274,274,274,274,274,274,274,257,1,1,274,274,274,274,1,0,1,257,1,1,1,1,257,257,1,1,1,1,1,1,257,274,274,274,274,274,274,274,274,274,274,530,546,546,819,1092,1365,1639,1912,2201,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2457,2168,1639,1365,1092,819,547,546,274,274,274,274,274,274,274,274,274,274,274,1,1,0,0,0,0,0,1,1,0,0,1,257,1,0,0,1,1,1,1,1,1,1,1,1,1,274,274,274,274,274,274,274,274,274,274,274,274,274,546,819,1092,1109,1639,1912,2185,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2458,2185,1911,1366,1093,819,547,546,274,274,274,257,1,1,1,257,257,257,257,1,1,0,0,0,0,0,0,0,1,0,0,0,274,1,0,0,1,1,1,1,1,1,1,1,1,1,257,1,1,1,1,1,257,257,257,1,274,274,274,274,546,819,820,1109,1639,1912,2201,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2459,2185,1912,1638,1349,820,547,546,274,274,274,274,257,1,1,1,1,257,257,1,1,1,0,0,0,0,0,0,0,274,0,0,0,274,1,0,0,1,1,1,1,1,1,1,1,1,1,257,1,1,1,1,1,1,274,1,1,1,274,274,274,274,546,547,836,1365,1639,1912,2185,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,4095,2457,2184,1639,1365,1092,803,530,274,274,274,274,274,257,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,257,274,0,0,0,1,1,1,0,1,1,1,1,1,257,1,1,1,1,257,1,1,1,0,1,1,274,1,0,1,274,274,274,274,274,274,563,836,1366,1639,1928,2184,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2441,2168,1639,1366,1093,820,547,274,274,257,257,257,1,1,1,1,1,1,1,1,1,1,1,0,256,256,0,0,0,1,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,1,1,1,1,1,1,1,1,1,1,1,1,1,274,274,274,274,274,546,563,1093,1366,1911,2185,2730,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2441,1912,1639,1366,1093,820,547,546,274,274,257,0,1,1,1,1,1,17,1,1,1,1,1,1,256,256,256,256,1,1,1,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,17,17,17,274,274,274,290,819,1109,1639,1912,2185,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2457,2168,1639,1366,1093,820,803,546,274,274,274,1,1,1,1,1,1,1,1,1,1,1,1,1,256,256,256,256,256,257,257,256,256,256,257,257,257,257,257,257,257,257,257,257,257,257,1,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,17,17,17,274,274,274,563,1092,1366,1639,1912,2185,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2457,2184,1895,1366,1093,820,803,546,274,274,274,274,274,1,1,1,1,1,1,1,1,0,0,0,256,256,256,256,256,256,256,256,272,272,274,274,274,274,274,274,274,257,257,257,257,257,256,256,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,17,274,274,274,547,820,1093,1366,1911,2184,2457,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,3003,2184,1895,1366,1093,820,547,546,274,274,274,274,274,17,1,1,1,0,0,0,0,0,256,256,256,256,272,274,274,529,529,529,529,529,529,529,529,529,529,529,529,529,529,529,529,274,257,256,257,257,257,257,1,1,1,1,1,1,1,1,1,0,0,0,0,0,1,1,274,274,274,546,819,1092,1365,1638,1911,2185,2457,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1895,1366,1092,819,547,546,274,274,274,257,257,1,1,0,0,0,0,0,0,256,256,272,272,274,529,529,529,529,529,801,801,801,801,801,801,801,801,801,801,801,801,801,785,785,529,529,529,529,274,274,257,257,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,274,274,274,546,819,1092,1365,1638,1912,2185,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1911,1366,1092,819,546,530,274,274,257,257,257,257,1,0,0,0,0,0,256,272,272,528,529,529,529,785,801,801,802,802,1058,1074,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1058,1058,1057,801,801,785,785,529,529,274,257,257,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,274,274,274,546,547,819,1092,1366,1639,1912,2201,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2457,1912,1639,1093,819,546,274,274,274,274,257,257,257,257,0,0,0,272,272,272,529,529,529,801,801,1057,1058,1058,1074,1330,1331,1331,1331,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1330,1330,1330,1330,1074,1058,1058,802,802,786,529,529,274,274,256,0,0,0,0,0,0,0,0,0,0,1,1,274,274,274,274,546,547,819,1093,1366,1639,2185,2730,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2459,2185,1911,1366,820,546,274,274,274,274,274,274,257,256,256,256,0,272,272,272,529,801,801,1057,1058,1330,1330,1330,1587,1603,1603,1603,1603,1859,1875,1875,1875,1859,1859,1859,1875,1875,1875,1859,1859,1859,1603,1603,1602,1586,1330,1330,1330,1058,1058,802,785,529,529,272,272,256,0,0,0,0,0,0,0,0,257,257,274,274,274,274,274,546,547,820,1093,1366,1912,2185,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,4095,2185,1912,1382,1093,819,546,274,274,274,274,274,274,274,272,272,274,274,529,545,801,801,1058,1074,1330,1330,1587,1603,1603,1859,1859,1860,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1875,1875,1859,1859,1859,1603,1603,1587,1331,1330,1330,1058,1058,801,801,529,529,272,256,0,0,0,0,256,256,256,256,257,274,274,274,274,274,274,547,820,1093,1638,1912,2185,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1912,1638,1093,820,547,546,274,274,274,272,272,274,274,274,274,529,545,801,801,1074,1330,1330,1603,1603,1859,1859,1859,1875,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2131,1875,1859,1859,1859,1859,1603,1603,1587,1330,1330,1074,801,801,529,272,256,256,256,256,256,257,256,256,257,274,274,257,274,274,274,290,547,820,1109,1639,2184,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2457,1912,1382,1109,820,563,546,274,274,272,272,272,272,529,529,529,529,801,1058,1074,1330,1331,1603,1603,1859,1876,1876,2132,2132,2132,2132,2132,2132,2132,2149,2148,2404,2404,2388,2388,2388,2388,2388,2404,2404,2404,2388,2388,2132,2132,2132,2132,2131,2131,2115,2115,1859,1859,1859,1603,1603,1330,1330,1058,801,801,529,529,256,256,257,256,256,256,256,257,257,257,1,1,274,274,290,819,1093,1366,1912,2185,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2457,2184,1639,1093,820,547,546,290,274,274,272,272,272,528,529,545,802,1058,1074,1331,1603,1603,1603,1876,1876,2132,2132,2132,2132,2132,2132,2132,2388,2388,2405,2405,2405,2405,2405,2404,2404,2404,2404,2404,2404,2404,2404,2404,2404,2388,2132,2132,2132,2132,2132,2132,2131,2131,2131,1859,1859,1859,1603,1603,1330,1330,1058,801,801,529,529,274,256,256,256,256,256,256,257,257,1,257,274,274,547,820,1093,1639,1928,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1639,1366,820,547,546,274,274,274,274,274,274,528,529,801,802,1074,1331,1603,1604,1876,1876,1876,2132,2132,2133,2133,2133,2133,2389,2389,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2404,2404,2404,2404,2404,2404,2388,2132,2132,2132,2132,2132,2132,2132,2131,2131,2131,1859,1859,1603,1603,1330,1330,1058,801,785,529,529,256,256,256,256,256,256,257,1,257,274,274,546,547,1092,1366,1912,2457,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1895,1366,1093,819,546,274,274,274,274,274,274,529,545,802,1074,1331,1347,1604,1876,1876,1876,2132,2133,2149,2149,2149,2149,2149,2133,2149,2149,2149,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2404,2404,2404,2404,2404,2404,2388,2388,2132,2132,2132,2132,2131,2131,2131,1875,1859,1859,1603,1603,1331,1074,1058,801,785,529,257,256,256,256,256,257,257,274,274,274,290,547,820,1109,1639,2185,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1912,1366,1093,820,546,274,274,274,274,274,274,529,801,802,1074,1331,1603,1876,1877,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2133,2149,2149,2149,2149,2149,2149,2149,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2404,2404,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1603,1587,1330,1058,801,785,529,257,256,256,256,257,257,274,274,274,274,290,563,1093,1366,1912,2187,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,4095,1912,1638,1093,819,547,530,530,274,274,274,274,529,545,802,1075,1347,1603,1876,1876,2133,2133,2149,2149,2149,2149,2133,2133,2133,2133,2133,2133,2133,2133,2149,2149,2149,2149,2149,2149,2149,2149,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2149,2148,2148,2148,2132,2132,2132,2132,2132,2132,2132,2132,2132,1860,1603,1603,1331,1330,1058,546,529,256,256,256,257,1,257,274,274,274,274,547,820,1366,1912,2458,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1639,1349,820,530,530,530,530,274,274,274,529,545,802,1075,1347,1604,1876,1876,2133,2149,2149,2133,2133,2133,2133,2133,1877,1877,1877,1877,1877,1877,1877,1877,1877,1893,2149,2149,2149,2149,2149,2149,2149,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2149,2149,2149,2149,2404,2388,2132,2132,2132,2132,2132,2132,2132,2132,1860,1859,1603,1603,1075,802,546,274,256,256,0,1,1,1,17,274,274,547,820,1093,1911,2441,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1912,1366,1092,803,274,530,530,530,530,530,529,529,802,802,1075,1348,1604,1620,1876,1876,1877,1876,1876,1876,1876,1876,1620,1604,1604,1604,1604,1604,1604,1604,1604,1620,1620,1620,1620,1877,1877,1893,2149,2149,2149,2149,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2149,2149,2149,2149,2149,2148,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1859,1859,1603,1331,1058,785,529,274,256,257,257,274,274,274,274,290,819,1093,1639,2185,2457,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,1912,1622,1349,819,546,274,274,274,530,530,530,546,546,803,1075,1075,1348,1348,1620,1620,1620,1620,1620,1604,1604,1348,1348,1347,1347,1331,1331,1331,1075,1075,1075,1075,1075,1347,1348,1348,1348,1604,1620,1877,1893,2149,2149,2149,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2149,2149,2149,2149,2149,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1603,1331,1058,801,529,274,274,274,274,274,274,274,274,547,1092,1638,2168,2457,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1638,1349,1076,803,546,274,530,530,530,546,546,803,803,819,1076,1348,1348,1604,1620,1621,1620,1620,1620,1348,1348,1348,1348,1348,1348,1331,1331,1075,1075,1075,1075,1075,1075,1075,1075,1075,1348,1348,1604,1620,1877,1877,2133,2133,2149,2149,2405,2405,2405,2405,2405,2405,2149,2149,2149,2149,2149,2149,2133,2133,2133,2132,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1860,1603,1331,1074,801,529,274,274,274,274,17,17,274,547,820,1365,1639,2184,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1911,1365,1076,803,546,546,546,546,547,547,547,803,803,819,1076,1348,1348,1605,1621,1877,1877,1877,1877,1621,1620,1620,1620,1604,1604,1604,1348,1348,1348,1348,1331,1331,1075,1075,1075,1075,1075,1075,1331,1348,1604,1604,1604,1877,1877,1877,2133,2133,2133,2149,2149,2149,2133,2133,2133,1877,1877,1877,1877,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,2132,2132,2133,2132,1876,1876,1860,1604,1331,1074,802,529,274,274,1,1,1,274,546,819,1092,1366,1911,2185,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1622,1092,803,546,530,546,546,547,803,803,803,803,819,1076,1092,1348,1605,1621,1877,1893,1893,1893,1877,1877,1877,1877,1877,1877,1621,1621,1621,1620,1604,1604,1348,1348,1347,1331,1331,1075,1075,1075,1331,1332,1332,1604,1604,1604,1604,1860,1877,1877,1877,1877,1877,1877,1877,1877,1877,1877,1621,1604,1604,1604,1604,1604,1604,1604,1604,1620,1620,1876,1876,1876,1877,1877,2133,2133,1877,1876,1876,1876,1604,1331,1074,546,529,274,1,1,1,274,274,547,819,1093,1638,1912,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1639,1349,819,546,530,274,530,546,547,803,803,803,819,1075,1076,1348,1349,1621,1877,1877,1893,1893,1893,1893,1893,1893,1893,1893,1893,1893,1893,1877,1877,1877,1877,1620,1604,1604,1348,1348,1347,1347,1332,1332,1332,1332,1332,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1348,1348,1348,1347,1331,1347,1347,1348,1348,1348,1604,1604,1604,1604,1620,1877,1877,1876,1876,1876,1877,1604,1348,1075,802,529,274,274,257,1,274,274,546,547,820,1366,1911,0,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1912,1366,1092,546,274,274,274,530,546,803,803,819,819,1075,1076,1348,1348,1621,1621,1877,1893,2150,2150,2149,2149,2149,2150,2150,2150,2150,2150,2150,2150,2150,2149,1893,1877,1877,1876,1604,1604,1604,1348,1604,1604,1588,1588,1332,1332,1332,1332,1332,1604,1604,1604,1604,1348,1348,1332,1332,1332,1332,1332,1331,1075,1075,1075,1075,1075,1075,1075,1075,1075,1331,1348,1348,1348,1348,1604,1604,1620,1876,1877,1877,1620,1604,1347,1075,802,529,274,274,1,274,274,274,290,547,1093,1639,2184,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1639,1093,819,546,274,274,274,529,546,802,819,819,1075,1076,1348,1348,1621,1621,1877,1893,1893,2150,2149,2149,2149,2149,2149,2150,2150,2150,2150,2150,2150,2150,2149,2149,2133,1877,1877,1876,1620,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1348,1347,1331,1331,1331,1332,1348,1348,1332,1332,1331,1331,1331,1348,1348,1348,1348,1348,1348,1348,1348,1348,1348,1604,1604,1620,1876,1876,1620,1604,1347,1075,818,802,529,274,274,274,274,274,274,547,1093,1382,1928,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,1912,1366,820,547,530,274,274,274,529,546,802,819,1075,1075,1348,1348,1605,1621,1877,1893,1894,2150,2149,2149,2149,2149,2149,2149,2149,2150,2406,2406,2406,2406,2150,2149,2149,2149,2133,1877,1877,1876,1876,1876,1876,1860,1860,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1347,1347,1331,1331,1331,1331,1348,1348,1348,1348,1348,1348,1348,1348,1348,1348,1348,1348,1348,1348,1348,1348,1348,1348,1604,1604,1604,1604,1604,1604,1348,1347,1075,802,546,529,274,274,17,17,274,291,820,1366,1912,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1639,1365,819,546,274,274,274,274,529,546,802,1075,1075,1348,1348,1621,1621,1877,1894,1894,2150,2150,2149,2149,2149,2149,2149,2149,2149,2405,2405,2406,2406,2149,2149,2149,2149,2149,2133,2133,1877,1876,1876,1876,1876,1876,1876,1860,1604,1604,1604,1604,1604,1604,1604,1604,1604,1603,1603,1331,1331,1331,1604,1604,1604,1604,1604,1604,1604,1620,1620,1620,1620,1620,1620,1620,1620,1604,1604,1604,1604,1604,1604,1620,1620,1620,1620,1604,1348,1075,1075,802,546,274,274,274,274,274,291,820,1109,1912,2730,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,1912,1366,1092,546,546,274,274,274,529,545,802,1075,1348,1348,1620,1621,1621,1877,1894,2150,2150,2150,2150,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2133,2133,2132,1876,1876,1876,1876,1876,1876,1876,1860,1860,1860,1860,1860,1876,1876,1876,1876,1860,1604,1603,1603,1603,1604,1604,1604,1876,1876,1877,1877,1877,1877,1877,1877,1877,1877,1877,1877,1877,1877,1877,1621,1621,1621,1620,1621,1877,1621,1620,1620,1348,1347,1075,802,546,546,274,274,274,274,290,820,1093,1655,2201,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,2457,1655,1109,819,546,274,274,274,529,545,802,1074,1347,1348,1620,1621,1877,1893,1894,2150,2150,2150,2150,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2133,2132,1876,1876,1876,1876,1876,1876,1876,1876,1876,1859,1859,1859,1860,1876,1876,1876,1876,1876,1876,1860,1603,1603,1604,1860,1860,1876,1876,1876,1877,1877,2133,2149,2149,2149,2149,2149,2149,2150,2149,2149,1893,1877,1877,1877,1877,1877,1877,1877,1877,1620,1604,1348,1075,818,802,546,546,546,290,290,291,820,1093,1639,2457,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,2185,1638,1092,819,274,274,274,529,545,801,1074,1347,1348,1620,1877,1893,1893,1893,2150,2150,2150,2150,2149,2149,1877,1877,1877,1877,1893,2149,2149,2149,2149,2149,2133,1877,1877,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1860,1603,1603,1859,1860,1876,2132,2132,2133,2132,1876,1860,1859,1587,1860,1860,1860,1876,1876,1876,1876,2133,2133,2149,2149,2149,2149,2149,2150,2150,2150,2150,2150,2149,1893,1893,1877,1877,1877,1877,1877,1621,1620,1348,1075,1075,819,803,803,547,547,547,547,820,1093,1639,2185,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,2184,1622,820,546,274,274,274,545,545,818,1075,1347,1620,1893,1893,1893,2149,2150,2150,2150,2150,2149,1893,1877,1877,1877,1877,1877,1877,1877,1876,1876,1876,1876,1876,1876,1876,1876,1620,1604,1604,1604,1860,1860,1876,1876,1876,1860,1860,1603,1603,1604,1860,1876,2133,2149,2149,2133,2132,1860,1859,1587,1860,1860,1860,1876,1876,1876,2132,2132,2133,2149,2149,2149,2149,2405,2406,2422,2422,2422,2150,2150,2150,2149,1893,1893,1893,1877,1877,1621,1620,1348,1348,1075,1075,819,819,820,820,820,820,1093,1365,1639,2185,4095,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,2457,1912,1365,819,546,274,529,529,545,818,1074,1347,1620,1876,1893,1893,2149,2149,2149,2149,2149,2149,2149,1877,1877,1876,1620,1620,1620,1620,1620,1604,1604,1604,1604,1604,1604,1604,1604,1603,1603,1603,1603,1604,1604,1604,1604,1604,1604,1603,1603,1603,1604,1860,2132,2149,2149,2405,2149,2132,1860,1859,1587,1604,1860,1860,1876,1876,1876,1876,2132,2132,2132,2149,2149,2149,2149,2406,2422,2422,2422,2150,2150,2150,2150,2149,1893,1877,1877,1877,1877,1621,1621,1348,1092,1076,1076,820,820,820,820,820,1092,1093,1639,2185,2458,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,2185,1639,1349,819,546,274,529,545,801,1074,1091,1347,1620,1893,2149,2149,2149,2149,1893,2149,2149,2149,1877,1877,1876,1604,1604,1604,1604,1604,1348,1347,1347,1331,1331,1331,1331,1331,1331,1331,1331,1331,1331,1331,1603,1604,1604,1604,1603,1587,1587,1587,1860,1876,2133,2405,2405,2405,2405,2132,1876,1603,1587,1604,1604,1860,1876,1876,1876,1876,1876,1876,2132,2132,2149,2149,2149,2406,2422,2422,2166,2166,2150,2150,2150,2149,1893,1877,1877,1877,1877,1621,1621,1349,1348,1092,1076,1076,820,820,820,820,1092,1093,1639,1912,2457,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,1912,1638,1092,803,546,274,529,545,802,1074,1347,1620,1876,1893,2149,2149,2149,2149,1893,1893,1893,2149,1877,1876,1620,1604,1604,1603,1347,1347,1331,1331,1331,1075,1075,1075,1075,1075,1075,1075,1075,1075,1331,1331,1348,1604,1604,1604,1603,1603,1603,1603,1860,2132,2149,2405,2405,2405,2405,2148,1876,1603,1331,1347,1604,1604,1604,1876,1876,1876,1876,1876,1876,1876,2132,2133,2149,2149,2150,2150,2150,2150,2150,2150,2150,2149,1893,1877,1877,1877,1877,1877,1621,1365,1348,1092,1076,1076,820,819,819,547,820,1092,1366,1639,2185,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,4095,1911,1365,820,546,545,274,529,545,818,1075,1347,1620,1892,2149,2165,2149,2149,1893,1893,1893,1893,1893,1877,1876,1604,1604,1347,1347,1331,1331,1075,1075,1075,1075,1075,1059,1075,1075,1075,1075,1075,1075,1075,1331,1332,1348,1604,1604,1604,1603,1603,1860,1876,2149,2405,2405,2405,2405,2405,2148,1876,1603,1331,1331,1331,1347,1604,1604,1604,1604,1604,1604,1860,1876,1876,1876,2133,2149,2149,2149,2149,2150,2150,2150,2149,2149,1893,1877,1893,1893,1894,1894,1621,1365,1348,1092,1076,819,819,803,547,546,547,820,1093,1366,1912,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,2457,1639,1093,819,546,529,529,545,801,818,1347,1603,1620,1892,2149,2149,2149,2149,2149,1893,1893,1893,2149,1877,1877,1876,1604,1604,1604,1347,1347,1331,1331,1075,1075,1075,1075,1075,1075,1075,1075,1075,1075,1331,1332,1348,1604,1605,1604,1604,1604,1860,1876,2133,2405,2405,2421,2421,2421,2405,2149,2148,1619,1347,1331,1331,1331,1603,1603,1603,1603,1603,1603,1603,1604,1604,1876,1876,1877,1877,1877,1893,1893,1893,1894,2149,2149,1893,1877,1893,1894,1894,1894,1621,1621,1349,1348,1076,819,819,547,546,274,546,547,1076,1366,1895,2730,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,2185,1638,1093,819,546,529,529,545,802,1074,1347,1620,1876,1893,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,1877,1877,1876,1620,1604,1604,1348,1348,1332,1331,1331,1331,1331,1331,1347,1348,1348,1348,1604,1604,1604,1877,1876,1620,1876,1876,1877,2149,2405,2405,2405,2421,2421,2405,2405,2149,1876,1603,1347,1331,1331,1347,1347,1331,1331,1331,1331,1331,1331,1348,1604,1604,1604,1621,1877,1877,1877,1877,1877,2149,2149,1877,1877,1893,1894,1894,1894,1878,1621,1621,1348,1348,1075,803,546,530,274,530,546,820,1349,1639,2184,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,2184,1622,1092,819,546,545,529,545,818,1090,1347,1620,1876,2149,2149,2149,2149,2149,2149,2149,2149,2149,2150,2150,2150,2150,2150,2149,1877,1877,1877,1620,1604,1604,1604,1604,1348,1348,1348,1604,1604,1604,1604,1604,1620,1876,1876,1877,1877,1876,1877,1877,2133,2405,2406,2405,2405,2405,2405,2405,2405,2405,2132,1859,1603,1331,1331,1331,1331,1331,1331,1075,1075,1075,1075,1331,1332,1348,1348,1604,1605,1605,1877,1877,1877,1877,1877,1877,1877,1877,1893,1894,1894,1893,1877,1621,1604,1348,1075,802,802,529,274,529,530,819,1093,1639,2185,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,0,1912,1366,1076,547,546,545,529,545,818,1090,1347,1620,1876,2149,2149,2149,2149,2149,2149,2149,2149,2150,2150,2150,2150,2150,2150,2149,2133,1877,1877,1877,1876,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1876,1876,1876,1876,1877,1877,2133,2133,2149,2405,2405,2405,2405,2405,2405,2405,2405,2405,2132,1876,1860,1603,1603,1603,1603,1331,1331,1331,1075,1075,1075,1075,1075,1075,1331,1332,1332,1348,1604,1604,1604,1877,1877,1877,1877,1877,1893,1894,1894,1894,1877,1877,1621,1348,1331,1075,802,545,529,530,546,819,1093,1638,2184,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,2186,1911,1365,820,547,546,545,545,801,818,1090,1347,1619,1876,2149,2149,2149,2149,2149,2149,2150,2150,2150,2406,2406,2406,2150,2149,2149,2133,1877,1877,1877,1877,1876,1876,1876,1860,1860,1604,1860,1860,1860,1876,1876,1876,1876,1876,1876,2132,2133,2149,2149,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2133,2132,1876,1860,1604,1603,1603,1331,1331,1331,1075,1075,1059,1059,1059,1059,1059,1059,1075,1331,1331,1331,1332,1604,1860,1876,1877,1877,1893,1893,1894,1894,1893,1877,1621,1604,1348,1075,802,802,545,546,802,819,1092,1638,2184,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,2185,1639,1093,819,546,546,545,545,802,1074,1091,1347,1620,1876,2149,2149,2149,2150,2406,2406,2406,2406,2406,2406,2406,2406,2406,2149,2149,2149,2133,2133,2133,2132,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,2132,2132,2132,2133,2133,2133,2149,2132,2132,2132,2132,2132,2132,2388,2388,2132,2132,2132,2132,2132,2132,1860,1860,1604,1604,1603,1347,1331,1331,1331,1075,1075,1075,1075,1075,1075,1075,1331,1331,1331,1332,1604,1604,1604,1604,1877,1877,1877,1893,1893,1877,1877,1621,1620,1348,1331,1074,802,801,802,803,1075,1092,1638,1928,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,2184,1638,1092,547,546,545,546,545,818,1074,1347,1363,1620,1893,2149,2150,2406,2422,2422,2422,2422,2422,2422,2406,2406,2406,2406,2405,2149,2149,2133,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2133,2149,2405,2149,2148,2132,2132,2132,2132,2116,2116,2132,2132,2132,2132,2132,2132,2132,2132,2132,2116,1860,1860,1604,1604,1604,1604,1347,1347,1331,1331,1331,1331,1075,1075,1331,1331,1331,1331,1331,1603,1603,1604,1604,1620,1877,1877,1877,1893,1877,1877,1877,1620,1604,1347,1075,1074,802,802,819,1075,1092,1366,1912,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,1912,1366,820,546,546,545,546,546,818,1091,1347,1620,1876,2149,2150,2406,2422,2422,2422,2422,2422,2422,2422,2406,2406,2406,2406,2405,2405,2405,2149,2149,2405,2405,2405,2405,2149,2149,2149,2149,2149,2149,2148,2132,2132,2132,2405,2405,2405,2132,2132,2132,2131,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,2116,2115,2115,1859,1860,1860,1604,1604,1604,1604,1604,1604,1348,1348,1348,1348,1331,1348,1604,1604,1604,1604,1604,1604,1604,1876,1876,1877,1877,1877,1893,1877,1877,1877,1876,1620,1347,1331,1074,802,818,819,1075,1092,1365,1911,2184,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,1912,1366,819,546,546,546,546,818,1075,1347,1620,1620,1893,2149,2422,2422,2422,2422,2422,2422,2422,2422,2422,2422,2406,2406,2406,2406,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2404,2404,2388,2388,2388,2388,2132,2131,1859,1858,1586,1586,1586,1586,1586,1587,1587,1587,1587,1587,1843,1859,1859,1859,1859,1859,1860,1860,1860,1860,1860,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1876,1877,1877,1877,1877,1877,1877,1893,1893,1893,1893,1893,1877,1877,1877,1620,1604,1347,1074,1074,1074,1075,1075,1092,1365,1911,2201,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,2184,1895,1365,819,546,546,546,546,818,1091,1348,1620,1893,2149,2150,2422,2422,2422,2422,2422,2422,2422,2422,2422,2422,2406,2406,2406,2406,2406,2405,2405,2405,2661,2661,2677,2677,2661,2405,2405,2405,2405,2405,2404,2404,2388,2388,2132,2132,2132,2131,1859,1586,1586,1313,1313,1313,1314,1330,1330,1586,1586,1586,1586,1586,1586,1843,1859,1859,1859,1860,1860,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1877,1877,1877,1877,2133,2149,2149,2149,2149,2149,2149,2149,2149,2149,1893,1877,1877,1876,1604,1347,1074,1074,1074,819,1075,1092,1365,1911,2185,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,2185,1639,1093,819,546,546,546,802,818,1091,1620,1620,1893,2165,2166,2422,2422,2422,2422,2422,2422,2422,2406,2406,2406,2406,2678,2678,2678,2678,2422,2422,2678,2677,2677,2677,2677,2677,2677,2405,2405,2405,2405,2404,2388,2132,2132,2132,2132,2131,1859,1586,1329,1313,1057,1057,1057,1313,1314,1314,1314,1314,1314,1314,1314,1314,1586,1859,1859,1859,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1877,1877,1877,2133,2133,2149,2150,2150,2150,2150,2150,2150,2149,2149,2149,2149,2133,1877,1876,1620,1347,1330,1074,1074,818,1075,1091,1365,1911,2185,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,2185,1639,1093,803,546,530,546,802,818,1347,1620,1893,2149,2166,2422,2422,2422,2422,2422,2422,2406,2406,2406,2406,2406,2406,2678,2678,2678,2678,2678,2678,2678,2678,2678,2678,2678,2677,2677,2405,2405,2405,2404,2388,2132,2132,2131,2115,2115,1859,1586,1329,1057,1040,784,1040,1041,1057,1057,1058,1058,1057,1057,1041,1057,1057,1314,1586,1859,1859,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,2132,2132,2133,2133,2133,2149,2149,2406,2406,2406,2406,2422,2422,2150,2150,2149,2149,2149,2149,2133,1876,1620,1603,1346,1074,1074,818,819,1075,1365,1655,2185,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,2185,1638,1093,803,546,530,546,802,1075,1348,1620,1893,2166,2166,2422,2422,2422,2422,2422,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2388,2132,2132,2132,1859,1859,1859,1859,1586,1313,1057,1040,1040,1057,1057,1057,1314,1058,1058,1057,1041,1041,1041,1041,1313,1586,1859,1859,2132,2132,2132,2132,2132,2132,2132,2132,2133,2133,2133,2133,2149,2149,2149,2149,2149,2149,2149,2406,2406,2406,2406,2406,2150,2149,2149,2149,2149,2133,1876,1620,1603,1347,1074,1074,818,818,819,1365,1655,2185,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,2185,1622,1092,803,546,530,546,802,1075,1348,1621,1893,2166,2422,2422,2422,2422,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2132,2132,2132,2116,1859,1859,1859,1586,1586,1330,1057,1057,1040,1040,1057,1314,1314,1314,1314,1058,1057,1041,785,784,784,1057,1330,1603,1859,2131,2132,2132,2132,2404,2404,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2149,2149,2133,2149,2149,2406,2406,2406,2406,2149,2149,2149,2149,2133,1876,1620,1603,1347,1330,1074,818,818,819,1092,1639,2184,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,2184,1366,1076,803,546,530,546,802,1075,1348,1877,2150,2166,2422,2422,2422,2422,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2388,2132,2132,2132,1859,1859,1859,1586,1586,1586,1329,1313,1057,1057,1313,1314,1330,1330,1330,1330,1314,1314,1057,1057,1041,784,1057,1330,1586,1859,2115,2131,2132,2132,2404,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2149,2405,2406,2406,2422,2422,2406,2406,2149,2149,2149,2149,1876,1620,1603,1347,1074,1074,818,818,819,1092,1638,2184,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,2168,1365,1076,546,530,530,546,802,1075,1348,1893,2150,2150,2166,2422,2422,2422,2406,2406,2406,2406,2406,2406,2406,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2132,2132,2132,2132,1859,1859,1859,1586,1586,1314,1313,1329,1330,1330,1330,1586,1587,1587,1587,1587,1587,1330,1314,1057,1057,1041,1057,1330,1586,1858,1859,2115,2131,2132,2404,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2406,2406,2422,2422,2422,2422,2150,2149,2149,2149,1876,1620,1603,1347,1074,1074,818,818,819,1092,1638,2184,273,273,273,273,273},
'{273,273,273,273,273,273,273,2184,1912,1349,819,546,530,546,546,819,1075,1604,1893,2150,2150,2150,2406,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2388,2132,2132,2132,2132,2115,1859,1859,1586,1586,1586,1586,1330,1586,1586,1587,1587,1587,1587,1587,1587,1587,1587,1330,1314,1313,1057,1313,1330,1586,1586,1859,1859,2131,2132,2404,2405,2405,2405,2405,2405,2405,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2422,2422,2422,2422,2406,2150,2149,2149,1876,1876,1603,1347,1074,1074,818,818,818,1092,1638,2184,273,273,273,273,273},
'{273,273,273,273,273,273,273,2730,1911,1093,819,546,530,546,802,819,1075,1620,1893,2150,2150,2150,2150,2149,2149,2149,2149,2149,2149,2405,2405,2405,2405,2405,2405,2405,2405,2149,2405,2405,2405,2405,2405,2405,2405,2404,2388,2132,2132,2132,2132,2132,2132,2115,1859,1859,1586,1586,1586,1586,1586,1587,1859,1859,1587,1587,1587,1587,1859,1859,1587,1586,1330,1313,1313,1330,1586,1586,1859,1859,2131,2132,2388,2405,2405,2405,2405,2405,2405,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2150,2149,2149,1877,1876,1603,1347,1074,1074,818,818,818,1092,1638,1928,273,273,273,273,273},
'{273,273,273,273,273,273,273,2441,1895,1092,819,546,530,546,802,1075,1348,1621,1894,2150,2150,2150,2149,2149,2149,2149,2149,2149,2149,2149,2405,2405,2405,2405,2405,2149,2149,2149,2149,2149,2149,2405,2148,2404,2388,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1859,1586,1586,1586,1843,1859,1859,1859,1843,1843,1843,1859,1859,1859,1859,1587,1586,1330,1330,1330,1586,1586,1859,1859,2132,2132,2132,2405,2405,2405,2405,2405,2405,2406,2406,2406,2406,2406,2406,2406,2422,2406,2406,2406,2406,2406,2406,2406,2406,2406,2149,2149,1893,1876,1620,1347,1074,1074,818,802,818,1092,1638,1928,273,273,273,273,273},
'{273,273,273,273,273,273,273,2458,1895,1092,803,546,530,530,802,1075,1348,1621,1894,2150,2150,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2405,2149,2149,2149,2149,2149,2149,2149,2149,2405,2405,2405,2405,2388,2132,2132,2132,2132,2132,2132,2132,2132,2132,2116,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1586,1586,1586,1586,1586,1859,1859,2115,2132,2132,2132,2405,2405,2405,2405,2405,2405,2405,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2149,2149,2149,2149,1876,1620,1347,1075,1074,802,802,802,1092,1382,1928,273,273,273,273,273},
'{273,273,273,273,273,273,273,2457,1639,1092,803,530,530,530,546,1075,1348,1621,1894,2150,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2133,2133,2133,2133,2133,2133,2133,2133,2405,2405,2405,2405,2404,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2116,2116,2116,2116,2116,2115,2115,2115,2115,2115,1859,1859,1859,1859,1843,1586,1586,1586,1586,1859,1859,2116,2132,2132,2132,2389,2405,2405,2405,2405,2405,2405,2405,2406,2405,2405,2405,2406,2406,2406,2406,2406,2406,2406,2422,2406,2405,2149,2149,2149,2149,1893,1876,1347,1331,1074,802,802,803,1092,1382,1912,273,273,273,273,273},
'{273,273,273,273,273,273,273,2457,1639,1092,803,530,530,530,802,1075,1348,1621,1894,2150,2149,2149,2149,2149,2133,2133,2133,2149,2133,2149,2149,2149,2133,2133,2133,2132,2132,2132,2132,2132,2132,2132,2132,2405,2405,2404,2388,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2116,2116,2115,2115,2115,2115,2115,2115,2115,2115,2115,2115,1859,1859,1859,1859,1859,1859,1859,1859,2116,2132,2132,2132,2132,2133,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2406,2406,2406,2406,2406,2406,2406,2406,2405,2149,2149,2149,2149,1893,1876,1604,1347,1074,802,802,802,1092,1382,1928,273,273,273,273,273},
'{273,273,273,273,273,273,273,2457,1639,1092,803,530,529,530,802,1075,1348,1621,1893,2150,2149,2149,2149,2133,2133,2132,2133,2133,2133,2133,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2404,2404,2388,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2116,2116,2115,2115,2115,2115,1843,1859,1859,1859,2115,2115,2115,2115,1859,1859,1859,1859,1859,2132,2132,2132,2132,2132,2133,2133,2133,2149,2149,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2406,2406,2406,2406,2149,2149,2149,2149,2149,1893,1877,1620,1347,1074,546,546,802,1092,1382,1928,273,273,273,273,273},
'{273,273,273,273,273,273,273,2457,1895,1092,819,546,529,546,802,1075,1348,1621,1893,1893,2149,2149,2149,2133,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2115,2115,1859,1859,1843,1843,1843,1843,1843,1843,1843,1843,1843,1843,1859,1859,1859,1859,1859,1859,1860,2116,2132,2132,2132,2132,2132,2389,2149,2149,2149,2149,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2149,2149,2405,2405,2149,2149,2149,2149,2149,2149,1877,1620,1347,1074,546,546,546,1092,1638,1928,273,273,273,273,273},
'{273,273,273,273,273,273,2971,2457,1895,1348,819,546,529,802,818,1075,1348,1621,1893,1893,2149,2149,2149,2149,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2116,2116,2115,1859,1859,1859,1842,1842,1842,1842,1842,1842,1842,1842,1842,1842,1842,1586,1842,1842,1843,1859,1859,2116,2132,2132,2132,2132,2132,2132,2132,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,1877,1620,1347,1074,545,546,546,1092,1638,2184,273,273,273,273,273},
'{273,273,273,273,273,273,2730,2441,1894,1348,1075,802,802,802,1075,1347,1620,1621,1877,1893,1893,2149,2149,2133,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2116,1859,1859,1859,1859,1859,1859,1843,1842,1586,1586,1570,1826,1826,1826,1826,1826,1826,1570,1570,1586,1586,1586,1842,1843,1859,1859,2116,2132,2132,2132,2132,2132,2132,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,1877,1620,1347,1074,529,546,802,1092,1638,2185,273,273,273,273,273},
'{273,273,273,273,273,2730,2713,2440,1894,1604,1347,1074,1074,1075,1347,1348,1620,1877,1893,1893,2149,2149,2149,2149,2148,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1859,1859,1859,1859,1843,1842,1842,1586,1586,1586,1842,1842,1842,1843,1842,1842,1842,1842,1842,1586,1586,1586,1586,1842,1843,1859,1859,1859,1860,2132,2132,2132,2132,2133,2405,2405,2405,2405,2405,2405,2405,2405,2149,2133,2133,2132,2132,2148,2149,2149,2149,2149,2149,2149,2149,2149,2133,2149,2149,2149,1893,1877,1604,1347,1074,529,546,547,1092,1639,2185,273,273,273,273,273},
'{273,273,273,273,0,2713,2440,2167,1894,1620,1348,1347,1347,1347,1604,1620,1876,1877,1893,2149,2149,2133,2149,2132,2148,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1843,1586,1586,1586,1586,1842,1586,1586,1586,1586,1842,1842,1843,1843,1843,1843,1843,1843,1842,1842,1842,1586,1586,1586,1586,1586,1586,1843,1859,1859,1859,2132,2132,2132,2132,2133,2405,2405,2405,2405,2405,2405,2149,2133,2132,2132,2132,2132,2132,2132,2132,2133,2133,2133,2133,2133,2133,2133,2133,2149,2149,1877,1877,1604,1347,802,529,546,803,1092,1639,2185,273,273,273,273,273},
'{273,273,273,273,2696,2423,2151,2150,1877,1604,1603,1603,1603,1604,1620,1876,1876,1877,1877,2133,2133,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1859,1586,1586,1586,1586,1586,1586,1842,1842,1842,1842,1843,1843,2115,2115,2115,2115,2099,1843,1843,1843,1843,1843,1842,1842,1842,1586,1586,1586,1587,1859,1859,1859,1860,2132,2132,2132,2133,2405,2405,2405,2405,2405,2149,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2133,2133,2133,2132,2132,2133,2133,1877,1877,1877,1604,1331,802,530,546,803,1093,1639,2185,273,273,273,273,273},
'{273,273,273,2696,2151,2133,1877,1860,1604,1603,1603,1876,1876,1876,1876,1876,1876,1877,2133,2133,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1586,1586,1586,1569,1570,1586,1586,1842,1843,1859,1859,2115,2115,2115,2115,2115,2115,2115,2115,2115,2115,2115,1859,1859,1859,1843,1586,1586,1586,1586,1587,1859,1859,1859,1859,2132,2132,2132,2132,2149,2149,2149,2405,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2133,1877,1877,1876,1604,1331,802,530,546,819,1093,1655,2186,273,273,273,273,273},
'{273,273,2696,2423,1877,1860,1603,1587,1587,1603,1603,1859,1860,1876,1876,1876,1876,1876,1877,1877,1877,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2131,1859,1859,1586,1586,1586,1586,1586,1586,1586,1843,1859,1859,1859,1859,1859,1859,1843,1843,1843,1843,1843,1843,1843,1843,1843,1843,1843,1843,1586,1586,1586,1586,1586,1586,1587,1603,1859,1859,1876,2132,2132,2149,2149,2149,2405,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1877,1877,1877,1620,1348,1331,802,530,546,819,1365,1911,2184,273,273,273,273,273},
'{273,2730,2423,2133,1860,1587,1570,1314,1586,1586,1603,1859,1859,1860,1876,1860,1860,1876,1876,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1859,1587,1586,1586,1586,1586,1843,1859,1859,1859,1859,1859,1859,1843,1842,1842,1842,1842,1586,1842,1842,1842,1842,1843,1843,1843,1587,1586,1586,1586,1586,1586,1586,1586,1586,1587,1859,1859,2132,2132,2132,2149,2149,2149,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1877,1877,1876,1604,1347,1075,802,530,803,820,1365,1912,0,273,273,273,273,273},
'{273,2423,2150,1860,1587,1570,1570,1570,1586,1586,1843,1859,1859,1859,1860,1860,1860,1876,1876,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1859,1859,1587,1843,1859,1859,1859,1859,1859,1859,1859,1859,1843,1842,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1314,1586,1586,1586,1603,1859,1876,2132,2132,2149,2149,2149,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1876,1876,1604,1331,1075,802,530,803,1076,1366,1912,273,273,273,273,273,273},
'{273,2423,1877,1859,1587,1586,1586,1586,1842,1842,1842,1859,1859,1859,1860,1860,1860,1876,1876,1876,1877,2132,2132,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1859,1859,1859,1859,1860,1860,1860,1860,1859,1859,1859,1587,1586,1586,1586,1586,1586,1586,1586,1570,1570,1570,1570,1570,1570,1586,1586,1586,1586,1586,1586,1586,1314,1586,1586,1586,1587,1859,1860,2132,2132,2149,2149,2149,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1876,1876,1876,1604,1331,1058,802,530,819,1092,1638,2185,273,273,273,273,273,273},
'{273,2150,1860,1843,1842,1842,1842,1842,1842,1843,1843,1843,1859,1859,1860,1860,1860,1876,1876,1876,1877,2132,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1860,1860,1876,2132,2132,1876,1860,1859,1859,1859,1587,1586,1586,1586,1586,1586,1586,1586,1570,1570,1570,1570,1570,1570,1586,1586,1586,1586,1587,1586,1586,1586,1586,1586,1586,1587,1859,1859,2132,2132,2132,2133,2149,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1876,1876,1604,1604,1331,1058,802,546,819,1349,1639,2185,273,273,273,273,273,273},
'{2184,2150,1860,1843,1842,1842,1842,2115,2115,2115,1859,1842,1859,1859,1860,1860,1860,1876,1876,1876,1876,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1860,1859,1859,1859,1859,1603,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1843,1843,1843,1859,1587,1587,1587,1587,1603,1603,1859,1859,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1876,1860,1604,1347,1075,1058,802,546,1076,1365,1911,2458,273,273,273,273,273,273},
'{2440,2150,1860,1843,1842,2098,2115,2115,2115,2115,1859,1842,1587,1859,1860,1860,1876,1620,1604,1876,1876,1876,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2131,2131,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1859,1859,1859,1859,1859,1859,1859,1587,1587,1586,1586,1586,1586,1586,1587,1843,1843,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,2132,1876,1876,1876,1876,1876,1860,1604,1331,1074,802,802,802,1076,1366,1912,2458,273,273,273,273,273,273},
'{2696,2406,1860,1843,1843,2099,2115,2115,2115,2115,1843,1586,1586,1603,1603,1860,1876,1876,1620,1876,1876,1876,1876,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1876,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1860,1860,1860,1859,1859,1859,1860,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1876,1876,1876,1860,1604,1331,1074,1058,802,802,1348,1638,2184,2457,273,273,273,273,273,273},
'{2680,2406,2116,1859,2115,2115,2115,2116,2115,1859,1842,1586,1586,1603,1603,1603,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1860,1860,1876,1876,2132,1876,1860,1859,1859,1859,1859,1859,1859,1859,1859,1860,2116,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1876,1876,1876,1604,1604,1347,1330,1058,1058,1075,1349,1895,2441,3983,273,273,273,273,273,273},
'{2696,2406,2133,2116,2115,2115,2115,2116,2115,1843,1586,1330,1330,1586,1603,1603,1604,1620,1620,1876,1876,1876,1876,1876,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1860,1860,1860,1860,1860,2116,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1860,1860,1876,1604,1604,1603,1331,1330,1331,1331,1621,1911,2440,2730,273,273,273,273,273,273},
'{2696,2406,2133,2116,2116,2115,2116,2116,1859,1842,1586,1313,1313,1330,1330,1603,1603,1604,1604,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1860,1860,1860,1860,1604,1604,1604,1603,1603,1603,1604,1877,2150,2440,2714,273,273,273,273,273,273},
'{2696,2422,2133,2132,2132,2115,2115,2115,1859,1586,1586,1313,1313,1330,1330,1587,1603,1604,1604,1860,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1860,1859,1603,1603,1603,1604,1604,1603,1603,1604,1604,1877,1894,2167,2440,273,273,273,273,273,273},
'{2696,2423,2405,2132,2132,2115,2115,2115,1842,1586,1313,1313,1313,1330,1330,1587,1603,1603,1860,1860,1860,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1860,1860,1860,1860,2116,2132,2132,1876,1876,2132,2132,2132,2132,2132,2132,2133,2133,2133,2133,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1859,1859,1603,1603,1603,1603,1603,1603,1603,1604,1604,1876,1877,2150,2167,2440,273,273,273,273,273},
'{2696,2423,2405,2132,2132,2115,2115,1859,1842,1586,1569,1313,1313,1330,1586,1587,1603,1603,1860,1860,1860,1876,1876,1876,1876,1876,1876,1876,1876,1875,1859,1859,1859,1859,1859,1859,1860,1860,2116,2132,1876,1876,2132,2132,2132,2132,2132,2133,2149,2405,2405,2405,2405,2149,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1860,1859,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1604,1876,1894,2167,2440,273,273,273,273},
'{2696,2423,2149,2132,2132,2115,2115,1858,1842,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1860,1860,1860,1860,1860,1860,1860,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1860,1860,1860,2132,1876,1876,2132,2132,2132,2132,2132,2148,2149,2405,2405,2405,2405,2405,2149,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1860,1860,1859,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1603,1587,1603,1876,1894,2423,273,273,273,273},
'{2696,2422,2149,2132,2132,2115,2115,1842,1842,1842,1842,1859,1859,1859,1859,1859,1603,1603,1603,1603,1604,1860,1860,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1860,1860,2116,2132,2132,2132,2132,2132,2132,2148,2148,2149,2405,2405,2405,2405,2405,2149,2148,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1860,1860,1860,1859,1859,1603,1603,1603,1603,1603,1603,1603,1858,1842,1586,1586,1586,1603,1876,2150,2730,273,273,273},
'{2440,2423,2149,2132,2132,2115,2115,2115,2115,1859,2115,2115,2115,2115,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1860,1860,1876,2132,2132,2132,2132,2132,2132,2148,2149,2149,2405,2405,2405,2405,2405,2149,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1860,1860,1860,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1858,1858,1842,1586,1586,1587,1860,2150,2440,273,273,273},
'{2184,2423,2149,2132,2132,2115,2115,2115,2115,2115,2132,2388,2132,2132,2132,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1860,1860,1876,2132,2132,2132,2132,2132,2132,2132,2149,2149,2405,2405,2405,2405,2405,2405,2132,2132,2132,2132,2132,2132,2132,1860,1859,1859,1859,2131,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,2132,2132,2132,2132,1876,1876,1876,1876,1876,1860,1860,1859,1859,1859,1603,1603,1603,1603,1603,1602,1602,1602,1603,1859,2114,1842,1842,1586,1587,1860,2150,2440,273,273,273},
'{273,2439,2150,2133,2132,2116,2115,2115,2116,2132,2132,2388,2132,2132,2132,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1860,1860,1876,2132,2132,2132,2132,2132,2132,2132,2132,2149,2149,2149,2405,2405,2149,2132,2132,2132,2132,2132,2132,1876,1860,1859,1859,1859,1859,1859,1875,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1876,1876,1876,1876,1860,1860,1860,1876,1860,1860,1859,1859,1603,1603,1603,1603,1587,1586,1586,1602,1603,1859,1859,2115,1859,1842,1843,1859,1860,2150,2424,273,273,273},
'{273,2440,2166,2149,2132,2116,2116,2116,2132,2132,2132,2132,2132,2115,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1860,1860,1860,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2149,2149,2149,2132,2132,2132,2132,2132,1876,1876,1860,1859,1859,1859,1859,1859,1859,1859,1859,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2131,1875,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1586,1586,1586,1586,1602,1603,1859,1859,2115,2115,1859,1859,1859,1860,2150,2424,273,273,273},
'{273,2184,2423,2150,2133,2132,2132,2132,2132,2132,2132,2116,1859,1859,1859,1603,1586,1586,1330,1347,1347,1347,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1860,1860,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1860,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1860,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2131,1875,1875,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1587,1586,1330,1586,1586,1586,1859,1859,2115,2115,2115,2115,1859,1860,1860,2150,2440,273,273,273},
'{273,273,2697,2423,2150,2133,2133,1876,1876,1860,1860,1859,1859,1587,1587,1586,1330,1330,1330,1330,1330,1331,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1876,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,1876,1876,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1860,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2131,1875,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1587,1586,1330,1330,1330,1586,1586,1603,1859,1859,2115,2116,2116,2116,1860,2133,2407,2696,273,273,273},
'{273,273,273,2440,2167,2150,2133,1877,1876,1860,1860,1603,1587,1587,1330,1330,1314,1330,1330,1330,1330,1330,1347,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1860,1876,1876,1876,1876,1876,1876,1876,1860,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1860,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2131,1875,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1587,1586,1330,1330,1330,1330,1586,1603,1859,1859,2116,2116,2116,2116,2116,2133,2423,2697,273,273,273},
'{273,273,273,273,2440,2423,2167,2150,1877,1877,1860,1604,1603,1587,1587,1330,1314,1314,1058,1330,1330,1331,1331,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1876,2132,2132,2132,2132,2132,2132,2131,1875,1875,1875,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1587,1587,1586,1330,1314,1314,1314,1330,1587,1859,1859,2116,2116,2116,2116,2133,2134,2424,2713,273,273,273},
'{273,273,273,273,273,2457,2440,2167,1894,1877,1877,1860,1604,1603,1587,1330,1314,1314,1058,1330,1331,1331,1331,1587,1587,1587,1587,1603,1603,1603,1586,1586,1586,1586,1586,1587,1587,1587,1587,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1587,1586,1586,1586,1586,1586,1586,1586,1586,1587,1587,1859,1859,1859,1859,1859,1859,1860,2132,1876,1875,1875,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1858,1858,1858,1602,1586,1586,1586,1587,1587,1587,1587,1330,1314,1314,1314,1330,1586,1603,1859,2116,2116,2116,2117,2133,2406,2440,273,273,273,273},
'{273,273,273,273,273,273,273,2440,2168,2167,1894,1894,1878,1877,1877,1348,1074,1058,1058,1074,1331,1331,1331,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1587,1587,1587,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1858,1858,1602,1602,1858,1858,1602,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1586,1586,1603,1859,2116,2116,2116,2133,2134,2407,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,2184,2184,2167,2167,1911,1621,1075,1075,1058,1074,1331,1331,1331,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1587,1587,1587,1587,1587,1587,1587,1587,1587,1587,1587,1587,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1602,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1858,1858,1586,1586,1586,1586,1858,1858,1586,1586,1586,1586,1586,1586,1330,1330,1330,1586,1587,1586,1586,1586,1586,1842,1859,2115,2116,2116,2133,2406,2440,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1638,1076,1075,1074,1074,1331,1331,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1587,1587,1587,1587,1587,1587,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1859,1859,1859,1859,1859,1602,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1586,1587,1587,1587,1842,1842,1843,1859,2115,2116,2116,2133,2406,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1894,1348,1075,1075,1075,1331,1331,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1330,1330,1314,1314,1314,1314,1314,1314,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1603,1603,1603,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1586,1587,1859,1859,1859,1859,1859,2115,2116,2116,2132,2149,2423,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1365,1092,1075,1075,1075,1331,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1313,1313,1314,1314,1314,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1586,1586,1859,1859,1859,2115,2115,2116,2116,2132,2133,2150,2423,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1638,1349,1075,1075,1075,1075,1331,1331,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1330,1330,1330,1314,1314,1314,1314,1314,1314,1058,1058,1058,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1313,1313,1313,1313,1314,1314,1314,1314,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1587,1859,1859,2115,2115,2116,2116,2133,2133,2150,2184,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1895,1365,1075,1075,1075,1075,1331,1347,1331,1330,1330,1330,1330,1330,1330,1330,1330,1074,1074,1074,1058,1058,1058,1314,1314,1314,1314,1314,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1058,1058,1057,1057,1313,1313,1313,1313,1314,1314,1314,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1330,1330,1330,1586,1586,1330,1330,1330,1330,1330,1330,1330,1074,1058,1058,1058,1330,1330,1330,1330,1586,1859,1859,2115,2132,2132,1860,1877,2133,2150,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1638,1092,1075,1075,1075,1331,1347,1331,1331,1331,1330,1330,1330,1330,1074,1074,1074,1074,1074,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1314,1314,1314,1314,1314,1314,1314,1314,1314,1058,1058,1058,1058,1058,1058,1058,1058,1058,1314,1058,1314,1314,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1074,1058,1058,1074,1331,1331,1603,1603,1603,1603,1859,1859,1860,1860,1876,1877,2150,2184,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1639,1349,1092,1076,1075,1347,1347,1331,1331,1331,1330,1330,1074,1074,1074,1074,1074,1074,1058,1058,1058,1058,1058,1058,1074,1074,1074,1074,1074,1074,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1314,1314,1314,1314,1314,1314,1314,1314,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1314,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1074,1058,1058,1058,1075,1331,1604,1604,1877,1604,1603,1587,1603,1860,1860,1877,1877,2150,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1911,1365,1348,1348,1348,1347,1347,1347,1331,1331,1331,1330,1074,1074,1074,1074,1074,1074,1074,1058,1058,1058,1058,1058,1074,1074,1074,1074,1074,1074,1074,1074,1058,1058,1058,1058,1058,1058,1058,1058,1314,1314,1314,1314,1314,1314,1314,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1074,1074,1074,1074,1075,1075,1348,1894,1894,2150,1894,1621,1604,1604,1860,1877,1894,2150,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1638,1365,1348,1348,1348,1347,1347,1331,1331,1331,1331,1331,1074,1074,1074,1074,1074,1074,1058,1058,1058,1058,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1058,1058,1058,1058,1058,1058,1058,1314,1314,1314,1314,1314,1314,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1074,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1074,1074,1075,1075,1075,1348,1622,2167,2440,2184,2168,1894,1878,1877,1877,1894,2167,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1895,1622,1349,1348,1348,1347,1347,1331,1331,1331,1331,1331,1331,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1058,1058,1058,1058,1058,1058,1314,1314,1314,1314,1314,1314,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1074,1330,1330,1330,1330,1074,1074,1074,1074,1074,1074,1074,1074,1074,1330,1074,1075,1075,1075,1075,1092,1365,1911,2184,273,273,273,273,2184,1895,1895,4095,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1641,1894,1621,1348,1348,1348,1347,1347,1331,1331,1331,1331,1331,1330,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1330,1074,1074,1074,1074,1074,1058,1058,1058,1058,1058,1314,1314,1314,1314,1314,1314,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1074,1074,1074,1075,1075,1075,1076,1349,1638,2457,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1911,1622,1349,1348,1348,1347,1347,1331,1331,1331,1331,1331,1330,1330,1330,1330,1074,1074,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1058,1058,1058,1314,1314,1314,1314,1314,1314,1314,1314,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1074,1074,1075,1075,1075,1092,1366,1912,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2168,1894,1621,1620,1604,1604,1603,1347,1331,1331,1331,1331,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1074,1075,1075,1092,1366,1911,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1895,1622,1621,1604,1604,1603,1603,1587,1331,1331,1331,1331,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1330,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1075,1092,1365,1639,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2168,1894,1877,1604,1604,1603,1603,1587,1587,1587,1331,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1330,1330,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1075,1075,1348,1638,2184,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1895,1877,1620,1604,1604,1603,1587,1587,1587,1587,1587,1587,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1314,1058,1058,1314,1314,1314,1314,1314,1314,1314,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1074,1075,1075,1075,1076,1365,1911,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2440,2167,1893,1876,1604,1604,1603,1603,1587,1587,1587,1587,1587,1587,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1330,1330,1330,1330,1314,1330,1330,1330,1330,1330,1330,1330,1314,1330,1074,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1074,1075,1075,1348,1348,1638,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2440,2167,1894,1876,1876,1604,1604,1603,1603,1603,1587,1587,1587,1587,1587,1587,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1330,1314,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1330,1074,1058,1058,1058,1058,1058,1058,1058,1058,1058,1074,1330,1075,1331,1348,1621,2409,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2730,2167,2150,1876,1876,1860,1604,1603,1603,1603,1603,1587,1587,1587,1587,1587,1331,1331,1331,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1314,1314,1314,1058,1058,1058,1314,1314,1314,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1058,1058,1058,1058,1058,1074,1330,1330,1330,1331,1331,1621,1894,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,2167,2150,1876,1876,1860,1604,1603,1603,1603,1603,1587,1587,1587,1587,1587,1587,1587,1331,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1074,1074,1074,1058,1074,1074,1330,1330,1331,1331,1348,1621,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,2150,1876,1876,1860,1604,1604,1603,1603,1603,1603,1587,1587,1587,1587,1587,1587,1587,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1314,1314,1314,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1074,1074,1074,1074,1330,1330,1331,1331,1347,1348,1622,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,2150,1876,1876,1860,1604,1603,1603,1603,1603,1603,1587,1587,1587,1587,1587,1587,1587,1587,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1074,1074,1074,1330,1330,1331,1331,1331,1347,1604,1894,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,2150,1876,1876,1860,1860,1603,1603,1603,1603,1603,1587,1587,1587,1587,1587,1587,1587,1587,1587,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1331,1331,1331,1347,1348,1620,1894,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,2150,1876,1876,1876,1860,1603,1603,1603,1603,1603,1603,1603,1587,1587,1587,1587,1587,1587,1587,1587,1587,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1331,1331,1331,1331,1347,1604,1621,1894,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,2149,1876,1876,1876,1860,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1587,1587,1587,1587,1587,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1331,1331,1331,1347,1603,1604,1621,1894,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,2149,1876,1876,1876,1860,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1587,1587,1587,1587,1587,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1331,1331,1331,1603,1603,1604,1621,1894,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,1893,1876,1876,1876,1860,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1587,1587,1587,1587,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1587,1603,1603,1603,1604,1621,1894,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,1893,1876,1876,1876,1860,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1587,1587,1587,1587,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1603,1603,1603,1603,1620,1621,1911,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2166,1893,1876,1876,1876,1860,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1587,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1620,1621,1911,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,2166,1893,1876,1876,1876,1860,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1602,1603,1603,1603,1603,1603,1620,1621,1911,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,4095,2166,1893,1876,1876,1876,1876,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1620,1621,1911,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2730,2150,1893,1876,1876,1876,1876,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1859,1603,1620,1637,1911,4095,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2457,2150,1893,1876,1876,1876,1876,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1603,1859,1603,1620,1637,1911,4095,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,2150,1893,1876,1876,1876,1876,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1587,1587,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1604,1620,1894,1911,2184,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,1894,1893,1876,1876,1876,1876,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1587,1603,1587,1587,1587,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1620,1620,1637,1911,1365,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,1894,1893,1876,1876,1876,1876,1859,1859,1859,1859,1859,1603,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1876,1620,1637,1911,2730,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,1894,1877,1876,1876,1876,1860,1859,1859,1859,1859,1859,1603,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1876,1620,1637,1911,1638,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,1894,1877,1876,1876,1876,1860,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1876,1876,1893,1910,2406,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1911,1894,1877,1876,1876,1876,1860,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1876,1876,1893,1910,2184,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1911,1894,1877,1876,1876,1876,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1876,1876,1893,1910,2167,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1911,1894,1877,1876,1876,1876,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1876,1876,1893,1894,2184,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,2167,1911,1894,1877,1876,1876,1860,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1876,1876,1877,1894,2168,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1912,1911,1911,1894,1894,1877,1876,1876,1860,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1876,1876,1877,1894,2168,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1656,1639,1639,1638,1894,1893,1877,1876,1876,1860,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1876,1876,1621,1894,2168,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1384,1367,1366,1366,1622,1621,1877,1876,1876,1876,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1876,1876,1621,1895,1912,273,273,273,273,273,273,273,273,273,2184,1657,1657,1657,1657,1657,1657,1641,1641,1384,1384,1385,1385,1641,1657,1657,1658},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,1384,1111,1093,1093,1093,1349,1621,1621,1876,1876,1876,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1876,1877,1621,1895,1912,1641,273,273,273,273,273,273,1657,1401,1385,1384,1384,1385,1385,1384,1384,1368,1368,1112,1112,1112,1112,1384,1385,1657,1658},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,1657,1111,1094,821,821,1092,1348,1621,1621,1876,1876,1876,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1860,1620,1621,1894,1896,1913,273,273,273,273,1675,1674,1402,1385,1385,1129,1112,1113,1113,1368,1368,1112,1112,1095,1095,1095,1112,1112,1385,1657,1658},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,1384,1094,821,548,820,1076,1348,1605,1620,1876,1876,1876,1859,1859,1875,1875,1875,1875,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1876,1620,1621,1622,1895,1912,1913,1930,1674,1675,1675,1659,1402,1385,1129,1113,1112,1113,1113,1112,1112,1096,839,839,839,839,839,1112,1385,1401,1658},
'{273,273,273,273,273,273,273,273,273,273,273,273,1913,1368,838,821,548,820,1076,1348,1604,1876,1876,1876,1876,1859,1859,1875,1875,1875,1875,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1860,1604,1621,1622,1639,1640,1657,1658,1658,1659,1659,1659,1402,1386,1385,1113,1113,1113,1113,1112,1112,840,839,839,839,839,840,1112,1385,1658,1931},
'{273,273,273,273,273,273,273,273,273,273,273,273,1657,1111,821,821,548,820,1348,1604,1620,1876,1876,1876,1876,1859,1859,1859,1859,1875,1875,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1587,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1587,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1604,1604,1621,1622,1639,1640,1641,1658,1658,1659,1659,1402,1402,1386,1129,1113,1113,1113,1112,1112,856,840,839,839,839,856,1113,1386,1658,1931},
'{273,273,273,273,273,273,273,273,273,273,273,4095,1640,1095,821,548,547,820,1348,1604,1876,1876,1876,1876,1876,1859,1859,1859,1859,1875,1875,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1587,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1604,1604,1621,1622,1623,1640,1641,1641,1658,1658,1659,1402,1402,1386,1129,1113,1113,1113,1113,1112,856,840,840,840,840,1112,1113,1402,1931,1948},
'{273,273,273,273,273,273,273,273,273,273,273,1914,1384,1094,549,548,547,1076,1348,1604,1876,1876,1876,1876,1875,1859,1859,1859,1859,1875,1875,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1876,1876,1876,1876,1859,1859,1859,1859,1859,1859,1604,1620,1621,1622,1367,1384,1385,1386,1402,1658,1402,1402,1386,1129,1113,1113,1113,1113,1113,857,856,840,840,840,1113,1385,1658,1931,2204},
'{273,273,273,273,273,273,273,273,273,273,273,1657,1367,822,548,548,547,1076,1348,1604,1876,1876,1876,1876,1875,1859,1859,1859,1859,1875,1875,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1876,1876,1876,1876,1876,1859,1859,1859,1859,1859,1859,1860,1620,1621,1622,1367,1367,1384,1385,1401,1658,1402,1386,1385,1113,1113,1113,1113,1113,1113,1113,857,856,856,856,1113,1386,1659,1932,2204},
'{273,273,273,273,273,273,273,273,273,273,273,1640,1367,821,548,804,803,1076,1604,1604,1876,1876,1876,1876,1875,1875,1875,1875,1875,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1876,1876,1876,1876,1876,1876,1875,1859,1859,1859,1859,1859,1860,1604,1621,1621,1622,1623,1639,1640,1641,1641,1641,1385,1385,1113,1112,1112,1112,1113,1113,1113,856,856,856,1113,1385,1658,1931,2204,2204},
'{273,273,273,273,273,273,273,273,273,273,2184,1384,1094,820,803,803,1076,1348,1604,1876,1876,1876,1876,1876,1876,1876,1875,1875,1875,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1586,1586,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1875,1876,1876,1876,1876,1876,1876,1876,1876,1859,1859,1859,1859,1859,1860,1860,1604,1621,1621,1622,1623,1623,1640,1640,1640,1624,1368,1368,1112,1112,1112,1112,1112,1112,856,1112,1113,1129,1386,1658,1931,2204,2204},
'{273,273,273,273,273,273,273,273,273,273,1929,1383,1094,820,803,1075,1332,1604,1604,1876,1876,1876,1876,1876,1876,1876,1875,1875,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1875,1876,1876,1876,1876,1876,1876,1876,1876,1859,1859,1859,1859,1859,1859,1860,1860,1621,1621,1622,1878,1879,1623,1623,1623,1368,1368,1367,1095,1095,839,840,1096,1096,840,1112,1113,1385,1402,1675,1931,2204,2204},
'{273,273,273,273,273,273,273,273,273,273,1657,1383,1094,1076,803,1075,1348,1604,1876,1876,1876,1876,1876,1875,1875,1875,1875,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1875,1876,1876,1876,1876,1876,1876,1876,1876,1859,1859,1859,1859,1859,1859,1859,1860,1860,1877,1877,1878,1878,1622,1623,1623,1367,1351,1095,1095,839,823,839,839,840,840,1096,1112,1385,1658,1931,1932,2204,2220},
'{273,273,273,273,273,273,273,273,273,273,1657,1367,1093,1076,1075,1331,1604,1604,1876,1876,1876,1876,1876,1875,1875,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1875,1876,1876,1876,1876,1876,1876,1876,1876,1859,1859,1859,1859,1859,1859,1859,1860,1860,1876,1877,1877,1877,1878,1622,1622,1606,1350,1094,1094,822,822,822,839,839,839,1096,1112,1385,1658,1931,1948,2204,2220},
'{273,273,273,273,273,273,273,273,273,273,1657,1367,1093,1076,1075,1347,1604,1876,1876,1876,1876,1876,1876,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1586,1586,1586,1586,1586,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1875,1876,1876,1876,1876,1876,1876,1876,1876,1859,1859,1859,1859,1859,1859,1859,1859,1860,1876,1876,1877,1877,1877,1877,1621,1605,1349,1349,1077,1077,821,822,822,823,1095,1096,1368,1385,1658,1931,1948,2204,2204}
};










parameter bit [11:0] HZColors2 [170][125] = '{
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,4095,2457,2457,2457,2457,2458,2458,2458,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2191,2459,2458,2185,2457,2457,2457,2185,2185,2184,1912,1912,2184,2184,2184,2185,2458,4095,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,2184,2184,2184,2185,2185,2185,2184,1912,1912,1912,1912,1912,1911,1639,1638,1638,1639,1639,1639,1911,2184,2185,2458,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2730,2457,2185,2184,1912,1639,1639,1639,1639,1911,1911,1639,1638,1638,1639,1638,1638,1366,1365,1093,1093,1365,1365,1365,1366,1639,1912,2185,2457,2458,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2186,2457,2185,2185,2184,1912,1911,1638,1366,1366,1366,1366,1366,1366,1366,1365,1365,1365,1365,1093,1093,1092,820,820,820,1092,1092,1093,1366,1639,1911,2184,2185,2185,2185,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2457,2185,2185,2185,2184,1912,1911,1911,1639,1638,1365,1093,1092,1092,1092,1092,1093,1092,820,820,820,820,820,820,819,547,547,547,547,547,819,1092,1365,1638,1911,1911,1912,1912,2185,2457,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2457,2185,2184,1912,1911,1639,1639,1638,1638,1366,1365,1365,1092,820,819,819,819,819,820,819,547,547,547,547,547,547,546,546,274,274,274,546,547,819,1092,1365,1638,1638,1638,1639,1912,2184,2457,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,2185,2184,1912,1911,1639,1638,1366,1365,1093,1093,1093,1092,1092,1092,819,547,547,546,546,547,547,546,546,546,546,546,546,546,530,274,274,274,274,274,546,547,819,1092,1365,1365,1365,1365,1638,1911,1912,2185,2457,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,2185,2184,1911,1639,1638,1366,1365,1093,820,820,819,819,819,819,819,819,547,546,530,274,274,274,530,274,274,274,274,274,274,274,274,274,274,274,274,274,274,546,547,819,1092,1092,820,1092,1093,1366,1639,1912,2184,2185,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1912,1911,1638,1366,1365,1093,1093,1092,820,819,547,546,546,546,546,546,546,546,274,274,274,274,274,274,274,274,274,274,274,274,274,274,274,274,274,274,274,274,274,546,547,819,819,819,819,820,1092,1365,1638,1639,1911,1912,2184,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1911,1638,1365,1093,1092,820,819,819,819,547,546,274,274,274,274,274,274,274,274,274,274,274,274,274,274,257,1,1,1,1,274,274,274,274,274,1,1,257,274,274,274,546,546,546,546,546,547,819,820,1093,1365,1365,1638,1911,1912,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1911,1638,1365,1092,820,819,547,547,547,546,546,274,274,274,274,274,274,274,274,274,274,274,274,274,274,257,1,1,1,1,1,274,274,274,274,257,1,1,1,274,274,274,274,274,274,274,274,530,546,547,820,820,1092,1093,1366,1638,1912,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1912,1638,1365,1092,819,547,546,546,274,274,530,274,274,274,274,274,274,274,274,274,274,274,274,274,274,1,1,1,257,1,1,1,257,274,274,274,1,1,1,1,1,274,274,274,274,274,274,274,274,274,546,546,547,547,819,1092,1365,1638,1912,2187,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1912,1638,1365,1092,819,547,546,274,274,274,274,274,274,274,274,274,274,274,274,257,1,1,274,274,274,274,1,0,1,257,1,1,1,1,257,257,1,1,1,1,1,1,257,274,274,274,274,274,274,274,274,274,274,530,546,546,819,1092,1365,1639,1912,2201,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2457,2168,1639,1365,1092,819,547,546,274,274,274,274,274,274,274,274,274,274,274,1,1,0,0,0,0,0,1,1,0,0,1,257,1,0,0,1,1,1,1,1,1,1,1,1,1,274,274,274,274,274,274,274,274,274,274,274,274,274,546,819,1092,1109,1639,1912,2185,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2458,2185,1911,1366,1093,819,547,546,274,274,274,257,1,1,1,257,257,257,257,1,1,0,0,0,0,0,0,0,1,0,0,0,274,1,0,0,1,1,1,1,1,1,1,1,1,1,257,1,1,1,1,1,257,257,257,1,274,274,274,274,546,819,820,1109,1639,1912,2201,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2459,2185,1912,1638,1349,820,547,546,274,274,274,274,257,1,1,1,1,257,257,1,1,1,0,0,0,0,0,0,0,274,0,0,0,274,1,0,0,1,1,1,1,1,1,1,1,1,1,257,1,1,1,1,1,1,274,1,1,1,274,274,274,274,546,547,836,1365,1639,1912,2185,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,4095,2457,2184,1639,1365,1092,803,530,274,274,274,274,274,257,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,257,274,0,0,0,1,1,1,0,1,1,1,1,1,257,1,1,1,1,257,1,1,1,0,1,1,274,1,0,1,274,274,274,274,274,274,563,836,1366,1639,1928,2184,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2441,2168,1639,1366,1093,820,547,274,274,257,257,257,1,1,1,1,1,1,1,1,1,1,1,0,256,256,0,0,0,1,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,1,1,1,1,1,1,1,1,1,1,1,1,1,274,274,274,274,274,546,563,1093,1366,1911,2185,2730,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2441,1912,1639,1366,1093,820,547,546,274,274,257,0,1,1,1,1,1,17,1,1,1,1,1,1,256,256,256,256,1,1,1,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,17,17,17,274,274,274,290,819,1109,1639,1912,2185,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2457,2168,1639,1366,1093,820,803,546,274,274,274,1,1,1,1,1,1,1,1,1,1,1,1,1,256,256,256,256,256,257,257,256,256,256,257,257,257,257,257,257,257,257,257,257,257,257,1,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,17,17,17,274,274,274,563,1092,1366,1639,1912,2185,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2457,2184,1895,1366,1093,820,803,546,274,274,274,274,274,1,1,1,1,1,1,1,1,0,0,0,256,256,256,256,256,256,256,256,272,272,274,274,274,274,274,274,274,257,257,257,257,257,256,256,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,17,274,274,274,547,820,1093,1366,1911,2184,2457,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,3003,2184,1895,1366,1093,820,547,546,274,274,274,274,274,17,1,1,1,0,0,0,0,0,256,256,256,256,272,274,274,529,529,529,529,529,529,529,529,529,529,529,529,529,529,529,529,274,257,256,257,257,257,257,1,1,1,1,1,1,1,1,1,0,0,0,0,0,1,1,274,274,274,546,819,1092,1365,1638,1911,2185,2457,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1895,1366,1092,819,547,546,274,274,274,257,257,1,1,0,0,0,0,0,0,256,256,272,272,274,529,529,529,529,529,801,801,801,801,801,801,801,801,801,801,801,801,801,785,785,529,529,529,529,274,274,257,257,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,274,274,274,546,819,1092,1365,1638,1912,2185,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1911,1366,1092,819,546,530,274,274,257,257,257,257,1,0,0,0,0,0,256,272,272,528,529,529,529,785,801,801,802,802,1058,1074,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1058,1058,1057,801,801,785,785,529,529,274,257,257,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,274,274,274,546,547,819,1092,1366,1639,1912,2201,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2457,1912,1639,1093,819,546,274,274,274,274,257,257,257,257,0,0,0,272,272,272,529,529,529,801,801,1057,1058,1058,1074,1330,1331,1331,1331,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1330,1330,1330,1330,1074,1058,1058,802,802,786,529,529,274,274,256,0,0,0,0,0,0,0,0,0,0,1,1,274,274,274,274,546,547,819,1093,1366,1639,2185,2730,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2459,2185,1911,1366,820,546,274,274,274,274,274,274,257,256,256,256,0,272,272,272,529,801,801,1057,1058,1330,1330,1330,1587,1603,1603,1603,1603,1859,1875,1875,1875,1859,1859,1859,1875,1875,1875,1859,1859,1859,1603,1603,1602,1586,1330,1330,1330,1058,1058,802,785,529,529,272,272,256,0,0,0,0,0,0,0,0,257,257,274,274,274,274,274,546,547,820,1093,1366,1912,2185,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,4095,2185,1912,1382,1093,819,546,274,274,274,274,274,274,274,272,272,274,274,529,545,801,801,1058,1074,1330,1330,1587,1603,1603,1859,1859,1860,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1875,1875,1859,1859,1859,1603,1603,1587,1331,1330,1330,1058,1058,801,801,529,529,272,256,0,0,0,0,256,256,256,256,257,274,274,274,274,274,274,547,820,1093,1638,1912,2185,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1912,1638,1093,820,547,546,274,274,274,272,272,274,274,274,274,529,545,801,801,1074,1330,1330,1603,1603,1859,1859,1859,1875,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2131,1875,1859,1859,1859,1859,1603,1603,1587,1330,1330,1074,801,801,529,272,256,256,256,256,256,257,256,256,257,274,274,257,274,274,274,290,547,820,1109,1639,2184,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2457,1912,1382,1109,820,563,546,274,274,272,272,272,272,529,529,529,529,801,1058,1074,1330,1331,1603,1603,1859,1876,1876,2132,2132,2132,2132,2132,2132,2132,2149,2148,2404,2404,2388,2388,2388,2388,2388,2404,2404,2404,2388,2388,2132,2132,2132,2132,2131,2131,2115,2115,1859,1859,1859,1603,1603,1330,1330,1058,801,801,529,529,256,256,257,256,256,256,256,257,257,257,1,1,274,274,290,819,1093,1366,1912,2185,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2457,2184,1639,1093,820,547,546,290,274,274,272,272,272,528,529,545,802,1058,1074,1331,1603,1603,1603,1876,1876,2132,2132,2132,2132,2132,2132,2132,2388,2388,2405,2405,2405,2405,2405,2404,2404,2404,2404,2404,2404,2404,2404,2404,2404,2388,2132,2132,2132,2132,2132,2132,2131,2131,2131,1859,1859,1859,1603,1603,1330,1330,1058,801,801,529,529,274,256,256,256,256,256,256,257,257,1,257,274,274,547,820,1093,1639,1928,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1639,1366,820,547,546,274,274,274,274,274,274,528,529,801,802,1074,1331,1603,1604,1876,1876,1876,2132,2132,2133,2133,2133,2133,2389,2389,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2404,2404,2404,2404,2404,2404,2388,2132,2132,2132,2132,2132,2132,2132,2131,2131,2131,1859,1859,1603,1603,1330,1330,1058,801,785,529,529,256,256,256,256,256,256,257,1,257,274,274,546,547,1092,1366,1912,2457,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1895,1366,1093,819,546,274,274,274,274,274,274,529,545,802,1074,1331,1347,1604,1876,1876,1876,2132,2133,2149,2149,2149,2149,2149,2133,2149,2149,2149,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2404,2404,2404,2404,2404,2404,2388,2388,2132,2132,2132,2132,2131,2131,2131,1875,1859,1859,1603,1603,1331,1074,1058,801,785,529,257,256,256,256,256,257,257,274,274,274,290,547,820,1109,1639,2185,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1912,1366,1093,820,546,274,274,274,274,274,274,529,801,802,1074,1331,1603,1876,1877,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2133,2149,2149,2149,2149,2149,2149,2149,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2404,2404,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1603,1587,1330,1058,801,785,529,257,256,256,256,257,257,274,274,274,274,290,563,1093,1366,1912,2187,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,4095,1912,1638,1093,819,547,530,530,274,274,274,274,529,545,802,1075,1347,1603,1876,1876,2133,2133,2149,2149,2149,2149,2133,2133,2133,2133,2133,2133,2133,2133,2149,2149,2149,2149,2149,2149,2149,2149,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2149,2148,2148,2148,2132,2132,2132,2132,2132,2132,2132,2132,2132,1860,1603,1603,1331,1330,1058,546,529,256,256,256,257,1,257,274,274,274,274,547,820,1366,1912,2458,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1639,1349,820,530,530,530,530,274,274,274,529,545,802,1075,1347,1604,1876,1876,2133,2149,2149,2133,2133,2133,2133,2133,1877,1877,1877,1877,1877,1877,1877,1877,1877,1893,2149,2149,2149,2149,2149,2149,2149,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2149,2149,2149,2149,2404,2388,2132,2132,2132,2132,2132,2132,2132,2132,1860,1859,1603,1603,1075,802,546,274,256,256,0,1,1,1,17,274,274,547,820,1093,1911,2441,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1912,1366,1092,803,274,530,530,530,530,530,529,529,802,802,1075,1348,1604,1620,1876,1876,1877,1876,1876,1876,1876,1876,1620,1604,1604,1604,1604,1604,1604,1604,1604,1620,1620,1620,1620,1877,1877,1893,2149,2149,2149,2149,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2149,2149,2149,2149,2149,2148,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1859,1859,1603,1331,1058,785,529,274,256,257,257,274,274,274,274,290,819,1093,1639,2185,2457,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,1912,1622,1349,819,546,274,274,274,530,530,530,546,546,803,1075,1075,1348,1348,1620,1620,1620,1620,1620,1604,1604,1348,1348,1347,1347,1331,1331,1331,1075,1075,1075,1075,1075,1347,1348,1348,1348,1604,1620,1877,1893,2149,2149,2149,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2149,2149,2149,2149,2149,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1603,1331,1058,801,529,274,274,274,274,274,274,274,274,547,1092,1638,2168,2457,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1638,1349,1076,803,546,274,530,530,530,546,546,803,803,819,1076,1348,1348,1604,1620,1621,1620,1620,1620,1348,1348,1348,1348,1348,1348,1331,1331,1075,1075,1075,1075,1075,1075,1075,1075,1075,1348,1348,1604,1620,1877,1877,2133,2133,2149,2149,2405,2405,2405,2405,2405,2405,2149,2149,2149,2149,2149,2149,2133,2133,2133,2132,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1860,1603,1331,1074,801,529,274,274,274,274,17,17,274,547,820,1365,1639,2184,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1911,1365,1076,803,546,546,546,546,547,547,547,803,803,819,1076,1348,1348,1605,1621,1877,1877,1877,1877,1621,1620,1620,1620,1604,1604,1604,1348,1348,1348,1348,1331,1331,1075,1075,1075,1075,1075,1075,1331,1348,1604,1604,1604,1877,1877,1877,2133,2133,2133,2149,2149,2149,2133,2133,2133,1877,1877,1877,1877,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,2132,2132,2133,2132,1876,1876,1860,1604,1331,1074,802,529,274,274,1,1,1,274,546,819,1092,1366,1911,2185,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1622,1092,803,546,530,546,546,547,803,803,803,803,819,1076,1092,1348,1605,1621,1877,1893,1893,1893,1877,1877,1877,1877,1877,1877,1621,1621,1621,1620,1604,1604,1348,1348,1347,1331,1331,1075,1075,1075,1331,1332,1332,1604,1604,1604,1604,1860,1877,1877,1877,1877,1877,1877,1877,1877,1877,1877,1621,1604,1604,1604,1604,1604,1604,1604,1604,1620,1620,1876,1876,1876,1877,1877,2133,2133,1877,1876,1876,1876,1604,1331,1074,546,529,274,1,1,1,274,274,547,819,1093,1638,1912,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1639,1349,819,546,530,274,530,546,547,803,803,803,819,1075,1076,1348,1349,1621,1877,1877,1893,1893,1893,1893,1893,1893,1893,1893,1893,1893,1893,1877,1877,1877,1877,1620,1604,1604,1348,1348,1347,1347,1332,1332,1332,1332,1332,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1348,1348,1348,1347,1331,1347,1347,1348,1348,1348,1604,1604,1604,1604,1620,1877,1877,1876,1876,1876,1877,1604,1348,1075,802,529,274,274,257,1,274,274,546,547,820,1366,1911,0,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1912,1366,1092,546,274,274,274,530,546,803,803,819,819,1075,1076,1348,1348,1621,1621,1877,1893,2150,2150,2149,2149,2149,2150,2150,2150,2150,2150,2150,2150,2150,2149,1893,1877,1877,1876,1604,1604,1604,1348,1604,1604,1588,1588,1332,1332,1332,1332,1332,1604,1604,1604,1604,1348,1348,1332,1332,1332,1332,1332,1331,1075,1075,1075,1075,1075,1075,1075,1075,1075,1331,1348,1348,1348,1348,1604,1604,1620,1876,1877,1877,1620,1604,1347,1075,802,529,274,274,1,274,274,274,290,547,1093,1639,2184,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1639,1093,819,546,274,274,274,529,546,802,819,819,1075,1076,1348,1348,1621,1621,1877,1893,1893,2150,2149,2149,2149,2149,2149,2150,2150,2150,2150,2150,2150,2150,2149,2149,2133,1877,1877,1876,1620,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1348,1347,1331,1331,1331,1332,1348,1348,1332,1332,1331,1331,1331,1348,1348,1348,1348,1348,1348,1348,1348,1348,1348,1604,1604,1620,1876,1876,1620,1604,1347,1075,818,802,529,274,274,274,274,274,274,547,1093,1382,1928,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,1912,1366,820,547,530,274,274,274,529,546,802,819,1075,1075,1348,1348,1605,1621,1877,1893,1894,2150,2149,2149,2149,2149,2149,2149,2149,2150,2406,2406,2406,2406,2150,2149,2149,2149,2133,1877,1877,1876,1876,1876,1876,1860,1860,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1347,1347,1331,1331,1331,1331,1348,1348,1348,1348,1348,1348,1348,1348,1348,1348,1348,1348,1348,1348,1348,1348,1348,1348,1604,1604,1604,1604,1604,1604,1348,1347,1075,802,546,529,274,274,17,17,274,291,820,1366,1912,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,2185,1639,1365,819,546,274,274,274,274,529,546,802,1075,1075,1348,1348,1621,1621,1877,1894,1894,2150,2150,2149,2149,2149,2149,2149,2149,2149,2405,2405,2406,2406,2149,2149,2149,2149,2149,2133,2133,1877,1876,1876,1876,1876,1876,1876,1860,1604,1604,1604,1604,1604,1604,1604,1604,1604,1603,1603,1331,1331,1331,1604,1604,1604,1604,1604,1604,1604,1620,1620,1620,1620,1620,1620,1620,1620,1604,1604,1604,1604,1604,1604,1620,1620,1620,1620,1604,1348,1075,1075,802,546,274,274,274,274,274,291,820,1109,1912,2730,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,1912,1366,1092,546,546,274,274,274,529,545,802,1075,1348,1348,1620,1621,1621,1877,1894,2150,2150,2150,2150,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2133,2133,2132,1876,1876,1876,1876,1876,1876,1876,1860,1860,1860,1860,1860,1876,1876,1876,1876,1860,1604,1603,1603,1603,1604,1604,1604,1876,1876,1877,1877,1877,1877,1877,1877,1877,1877,1877,1877,1877,1877,1877,1621,1621,1621,1620,1621,1877,1621,1620,1620,1348,1347,1075,802,546,546,274,274,274,274,290,820,1093,1655,2201,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,2457,1655,1109,819,546,274,274,274,529,545,802,1074,1347,1348,1620,1621,1877,1893,1894,2150,2150,2150,2150,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2133,2132,1876,1876,1876,1876,1876,1876,1876,1876,1876,1859,1859,1859,1860,1876,1876,1876,1876,1876,1876,1860,1603,1603,1604,1860,1860,1876,1876,1876,1877,1877,2133,2149,2149,2149,2149,2149,2149,2150,2149,2149,1893,1877,1877,1877,1877,1877,1877,1877,1877,1620,1604,1348,1075,818,802,546,546,546,290,290,291,820,1093,1639,2457,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,2185,1638,1092,819,274,274,274,529,545,801,1074,1347,1348,1620,1877,1893,1893,1893,2150,2150,2150,2150,2149,2149,1877,1877,1877,1877,1893,2149,2149,2149,2149,2149,2133,1877,1877,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1860,1603,1603,1859,1860,1876,2132,2132,2133,2132,1876,1860,1859,1587,1860,1860,1860,1876,1876,1876,1876,2133,2133,2149,2149,2149,2149,2149,2150,2150,2150,2150,2150,2149,1893,1893,1877,1877,1877,1877,1877,1621,1620,1348,1075,1075,819,803,803,547,547,547,547,820,1093,1639,2185,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,2184,1622,820,546,274,274,274,545,545,818,1075,1347,1620,1893,1893,1893,2149,2150,2150,2150,2150,2149,1893,1877,1877,1877,1877,1877,1877,1877,1876,1876,1876,1876,1876,1876,1876,1876,1620,1604,1604,1604,1860,1860,1876,1876,1876,1860,1860,1603,1603,1604,1860,1876,2133,2149,2149,2133,2132,1860,1859,1587,1860,1860,1860,1876,1876,1876,2132,2132,2133,2149,2149,2149,2149,2405,2406,2422,2422,2422,2150,2150,2150,2149,1893,1893,1893,1877,1877,1621,1620,1348,1348,1075,1075,819,819,820,820,820,820,1093,1365,1639,2185,4095,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,2457,1912,1365,819,546,274,529,529,545,818,1074,1347,1620,1876,1893,1893,2149,2149,2149,2149,2149,2149,2149,1877,1877,1876,1620,1620,1620,1620,1620,1604,1604,1604,1604,1604,1604,1604,1604,1603,1603,1603,1603,1604,1604,1604,1604,1604,1604,1603,1603,1603,1604,1860,2132,2149,2149,2405,2149,2132,1860,1859,1587,1604,1860,1860,1876,1876,1876,1876,2132,2132,2132,2149,2149,2149,2149,2406,2422,2422,2422,2150,2150,2150,2150,2149,1893,1877,1877,1877,1877,1621,1621,1348,1092,1076,1076,820,820,820,820,820,1092,1093,1639,2185,2458,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,2185,1639,1349,819,546,274,529,545,801,1074,1091,1347,1620,1893,2149,2149,2149,2149,1893,2149,2149,2149,1877,1877,1876,1604,1604,1604,1604,1604,1348,1347,1347,1331,1331,1331,1331,1331,1331,1331,1331,1331,1331,1331,1603,1604,1604,1604,1603,1587,1587,1587,1860,1876,2133,2405,2405,2405,2405,2132,1876,1603,1587,1604,1604,1860,1876,1876,1876,1876,1876,1876,2132,2132,2149,2149,2149,2406,2422,2422,2166,2166,2150,2150,2150,2149,1893,1877,1877,1877,1877,1621,1621,1349,1348,1092,1076,1076,820,820,820,820,1092,1093,1639,1912,2457,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,1912,1638,1092,803,546,274,529,545,802,1074,1347,1620,1876,1893,2149,2149,2149,2149,1893,1893,1893,2149,1877,1876,1620,1604,1604,1603,1347,1347,1331,1331,1331,1075,1075,1075,1075,1075,1075,1075,1075,1075,1331,1331,1348,1604,1604,1604,1603,1603,1603,1603,1860,2132,2149,2405,2405,2405,2405,2148,1876,1603,1331,1347,1604,1604,1604,1876,1876,1876,1876,1876,1876,1876,2132,2133,2149,2149,2150,2150,2150,2150,2150,2150,2150,2149,1893,1877,1877,1877,1877,1877,1621,1365,1348,1092,1076,1076,820,819,819,547,820,1092,1366,1639,2185,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,4095,1911,1365,820,546,545,274,529,545,818,1075,1347,1620,1892,2149,2165,2149,2149,1893,1893,1893,1893,1893,1877,1876,1604,1604,1347,1347,1331,1331,1075,1075,1075,1075,1075,1059,1075,1075,1075,1075,1075,1075,1075,1331,1332,1348,1604,1604,1604,1603,1603,1860,1876,2149,2405,2405,2405,2405,2405,2148,1876,1603,1331,1331,1331,1347,1604,1604,1604,1604,1604,1604,1860,1876,1876,1876,2133,2149,2149,2149,2149,2150,2150,2150,2149,2149,1893,1877,1893,1893,1894,1894,1621,1365,1348,1092,1076,819,819,803,547,546,547,820,1093,1366,1912,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,2457,1639,1093,819,546,529,529,545,801,818,1347,1603,1620,1892,2149,2149,2149,2149,2149,1893,1893,1893,2149,1877,1877,1876,1604,1604,1604,1347,1347,1331,1331,1075,1075,1075,1075,1075,1075,1075,1075,1075,1075,1331,1332,1348,1604,1605,1604,1604,1604,1860,1876,2133,2405,2405,2421,2421,2421,2405,2149,2148,1619,1347,1331,1331,1331,1603,1603,1603,1603,1603,1603,1603,1604,1604,1876,1876,1877,1877,1877,1893,1893,1893,1894,2149,2149,1893,1877,1893,1894,1894,1894,1621,1621,1349,1348,1076,819,819,547,546,274,546,547,1076,1366,1895,2730,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,2185,1638,1093,819,546,529,529,545,802,1074,1347,1620,1876,1893,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,1877,1877,1876,1620,1604,1604,1348,1348,1332,1331,1331,1331,1331,1331,1347,1348,1348,1348,1604,1604,1604,1877,1876,1620,1876,1876,1877,2149,2405,2405,2405,2421,2421,2405,2405,2149,1876,1603,1347,1331,1331,1347,1347,1331,1331,1331,1331,1331,1331,1348,1604,1604,1604,1621,1877,1877,1877,1877,1877,2149,2149,1877,1877,1893,1894,1894,1894,1878,1621,1621,1348,1348,1075,803,546,530,274,530,546,820,1349,1639,2184,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,2184,1622,1092,819,546,545,529,545,818,1090,1347,1620,1876,2149,2149,2149,2149,2149,2149,2149,2149,2149,2150,2150,2150,2150,2150,2149,1877,1877,1877,1620,1604,1604,1604,1604,1348,1348,1348,1604,1604,1604,1604,1604,1620,1876,1876,1877,1877,1876,1877,1877,2133,2405,2406,2405,2405,2405,2405,2405,2405,2405,2132,1859,1603,1331,1331,1331,1331,1331,1331,1075,1075,1075,1075,1331,1332,1348,1348,1604,1605,1605,1877,1877,1877,1877,1877,1877,1877,1877,1893,1894,1894,1893,1877,1621,1604,1348,1075,802,802,529,274,529,530,819,1093,1639,2185,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,0,1912,1366,1076,547,546,545,529,545,818,1090,1347,1620,1876,2149,2149,2149,2149,2149,2149,2149,2149,2150,2150,2150,2150,2150,2150,2149,2133,1877,1877,1877,1876,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1876,1876,1876,1876,1877,1877,2133,2133,2149,2405,2405,2405,2405,2405,2405,2405,2405,2405,2132,1876,1860,1603,1603,1603,1603,1331,1331,1331,1075,1075,1075,1075,1075,1075,1331,1332,1332,1348,1604,1604,1604,1877,1877,1877,1877,1877,1893,1894,1894,1894,1877,1877,1621,1348,1331,1075,802,545,529,530,546,819,1093,1638,2184,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,2186,1911,1365,820,547,546,545,545,801,818,1090,1347,1619,1876,2149,2149,2149,2149,2149,2149,2150,2150,2150,2406,2406,2406,2150,2149,2149,2133,1877,1877,1877,1877,1876,1876,1876,1860,1860,1604,1860,1860,1860,1876,1876,1876,1876,1876,1876,2132,2133,2149,2149,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2133,2132,1876,1860,1604,1603,1603,1331,1331,1331,1075,1075,1059,1059,1059,1059,1059,1059,1075,1331,1331,1331,1332,1604,1860,1876,1877,1877,1893,1893,1894,1894,1893,1877,1621,1604,1348,1075,802,802,545,546,802,819,1092,1638,2184,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,2185,1639,1093,819,546,546,545,545,802,1074,1091,1347,1620,1876,2149,2149,2149,2150,2406,2406,2406,2406,2406,2406,2406,2406,2406,2149,2149,2149,2133,2133,2133,2132,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,2132,2132,2132,2133,2133,2133,2149,2132,2132,2132,2132,2132,2132,2388,2388,2132,2132,2132,2132,2132,2132,1860,1860,1604,1604,1603,1347,1331,1331,1331,1075,1075,1075,1075,1075,1075,1075,1331,1331,1331,1332,1604,1604,1604,1604,1877,1877,1877,1893,1893,1877,1877,1621,1620,1348,1331,1074,802,801,802,803,1075,1092,1638,1928,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,2184,1638,1092,547,546,545,546,545,818,1074,1347,1363,1620,1893,2149,2150,2406,2422,2422,2422,2422,2422,2422,2406,2406,2406,2406,2405,2149,2149,2133,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2133,2149,2405,2149,2148,2132,2132,2132,2132,2116,2116,2132,2132,2132,2132,2132,2132,2132,2132,2132,2116,1860,1860,1604,1604,1604,1604,1347,1347,1331,1331,1331,1331,1075,1075,1331,1331,1331,1331,1331,1603,1603,1604,1604,1620,1877,1877,1877,1893,1877,1877,1877,1620,1604,1347,1075,1074,802,802,819,1075,1092,1366,1912,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,1912,1366,820,546,546,545,546,546,818,1091,1347,1620,1876,2149,2150,2406,2422,2422,2422,2422,2422,2422,2422,2406,2406,2406,2406,2405,2405,2405,2149,2149,2405,2405,2405,2405,2149,2149,2149,2149,2149,2149,2148,2132,2132,2132,2405,2405,2405,2132,2132,2132,2131,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,2116,2115,2115,1859,1860,1860,1604,1604,1604,1604,1604,1604,1348,1348,1348,1348,1331,1348,1604,1604,1604,1604,1604,1604,1604,1876,1876,1877,1877,1877,1893,1877,1877,1877,1876,1620,1347,1331,1074,802,818,819,1075,1092,1365,1911,2184,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,1912,1366,819,546,546,546,546,818,1075,1347,1620,1620,1893,2149,2422,2422,2422,2422,2422,2422,2422,2422,2422,2422,2406,2406,2406,2406,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2404,2404,2388,2388,2388,2388,2132,2131,1859,1858,1586,1586,1586,1586,1586,1587,1587,1587,1587,1587,1843,1859,1859,1859,1859,1859,1860,1860,1860,1860,1860,1604,1604,1604,1604,1604,1604,1604,1604,1604,1604,1876,1877,1877,1877,1877,1877,1877,1893,1893,1893,1893,1893,1877,1877,1877,1620,1604,1347,1074,1074,1074,1075,1075,1092,1365,1911,2201,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,2184,1895,1365,819,546,546,546,546,818,1091,1348,1620,1893,2149,2150,2422,2422,2422,2422,2422,2422,2422,2422,2422,2422,2406,2406,2406,2406,2406,2405,2405,2405,2661,2661,2677,2677,2661,2405,2405,2405,2405,2405,2404,2404,2388,2388,2132,2132,2132,2131,1859,1586,1586,1313,1313,1313,1314,1330,1330,1586,1586,1586,1586,1586,1586,1843,1859,1859,1859,1860,1860,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1877,1877,1877,1877,2133,2149,2149,2149,2149,2149,2149,2149,2149,2149,1893,1877,1877,1876,1604,1347,1074,1074,1074,819,1075,1092,1365,1911,2185,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,2185,1639,1093,819,546,546,546,802,818,1091,1620,1620,1893,2165,2166,2422,2422,2422,2422,2422,2422,2422,2406,2406,2406,2406,2678,2678,2678,2678,2422,2422,2678,2677,2677,2677,2677,2677,2677,2405,2405,2405,2405,2404,2388,2132,2132,2132,2132,2131,1859,1586,1329,1313,1057,1057,1057,1313,1314,1314,1314,1314,1314,1314,1314,1314,1586,1859,1859,1859,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1877,1877,1877,2133,2133,2149,2150,2150,2150,2150,2150,2150,2149,2149,2149,2149,2133,1877,1876,1620,1347,1330,1074,1074,818,1075,1091,1365,1911,2185,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,2185,1639,1093,803,546,530,546,802,818,1347,1620,1893,2149,2166,2422,2422,2422,2422,2422,2422,2406,2406,2406,2406,2406,2406,2678,2678,2678,2678,2678,2678,2678,2678,2678,2678,2678,2677,2677,2405,2405,2405,2404,2388,2132,2132,2131,2115,2115,1859,1586,1329,1057,1040,784,1040,1041,1057,1057,1058,1058,1057,1057,1041,1057,1057,1314,1586,1859,1859,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,2132,2132,2133,2133,2133,2149,2149,2406,2406,2406,2406,2422,2422,2150,2150,2149,2149,2149,2149,2133,1876,1620,1603,1346,1074,1074,818,819,1075,1365,1655,2185,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,2185,1638,1093,803,546,530,546,802,1075,1348,1620,1893,2166,2166,2422,2422,2422,2422,2422,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2388,2132,2132,2132,1859,1859,1859,1859,1586,1313,1057,1040,1040,1057,1057,1057,1314,1058,1058,1057,1041,1041,1041,1041,1313,1586,1859,1859,2132,2132,2132,2132,2132,2132,2132,2132,2133,2133,2133,2133,2149,2149,2149,2149,2149,2149,2149,2406,2406,2406,2406,2406,2150,2149,2149,2149,2149,2133,1876,1620,1603,1347,1074,1074,818,818,819,1365,1655,2185,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,2185,1622,1092,803,546,530,546,802,1075,1348,1621,1893,2166,2422,2422,2422,2422,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2132,2132,2132,2116,1859,1859,1859,1586,1586,1330,1057,1057,1040,1040,1057,1314,1314,1314,1314,1058,1057,1041,785,784,784,1057,1330,1603,1859,2131,2132,2132,2132,2404,2404,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2149,2149,2133,2149,2149,2406,2406,2406,2406,2149,2149,2149,2149,2133,1876,1620,1603,1347,1330,1074,818,818,819,1092,1639,2184,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,2184,1366,1076,803,546,530,546,802,1075,1348,1877,2150,2166,2422,2422,2422,2422,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2388,2132,2132,2132,1859,1859,1859,1586,1586,1586,1329,1313,1057,1057,1313,1314,1330,1330,1330,1330,1314,1314,1057,1057,1041,784,1057,1330,1586,1859,2115,2131,2132,2132,2404,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2149,2405,2406,2406,2422,2422,2406,2406,2149,2149,2149,2149,1876,1620,1603,1347,1074,1074,818,818,819,1092,1638,2184,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,2168,1365,1076,546,530,530,546,802,1075,1348,1893,2150,2150,2166,2422,2422,2422,2406,2406,2406,2406,2406,2406,2406,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2132,2132,2132,2132,1859,1859,1859,1586,1586,1314,1313,1329,1330,1330,1330,1586,1587,1587,1587,1587,1587,1330,1314,1057,1057,1041,1057,1330,1586,1858,1859,2115,2131,2132,2404,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2406,2406,2422,2422,2422,2422,2150,2149,2149,2149,1876,1620,1603,1347,1074,1074,818,818,819,1092,1638,2184,273,273,273,273,273},
'{273,273,273,273,273,273,273,2184,1912,1349,819,546,530,546,546,819,1075,1604,1893,2150,2150,2150,2406,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2388,2132,2132,2132,2132,2115,1859,1859,1586,1586,1586,1586,1330,1586,1586,1587,1587,1587,1587,1587,1587,1587,1587,1330,1314,1313,1057,1313,1330,1586,1586,1859,1859,2131,2132,2404,2405,2405,2405,2405,2405,2405,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2422,2422,2422,2422,2406,2150,2149,2149,1876,1876,1603,1347,1074,1074,818,818,818,1092,1638,2184,273,273,273,273,273},
'{273,273,273,273,273,273,273,2730,1911,1093,819,546,530,546,802,819,1075,1620,1893,2150,2150,2150,2150,2149,2149,2149,2149,2149,2149,2405,2405,2405,2405,2405,2405,2405,2405,2149,2405,2405,2405,2405,2405,2405,2405,2404,2388,2132,2132,2132,2132,2132,2132,2115,1859,1859,1586,1586,1586,1586,1586,1587,1859,1859,1587,1587,1587,1587,1859,1859,1587,1586,1330,1313,1313,1330,1586,1586,1859,1859,2131,2132,2388,2405,2405,2405,2405,2405,2405,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2150,2149,2149,1877,1876,1603,1347,1074,1074,818,818,818,1092,1638,1928,273,273,273,273,273},
'{273,273,273,273,273,273,273,2441,1895,1092,819,546,530,546,802,1075,1348,1621,1894,2150,2150,2150,2149,2149,2149,2149,2149,2149,2149,2149,2405,2405,2405,2405,2405,2149,2149,2149,2149,2149,2149,2405,2148,2404,2388,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1859,1586,1586,1586,1843,1859,1859,1859,1843,1843,1843,1859,1859,1859,1859,1587,1586,1330,1330,1330,1586,1586,1859,1859,2132,2132,2132,2405,2405,2405,2405,2405,2405,2406,2406,2406,2406,2406,2406,2406,2422,2406,2406,2406,2406,2406,2406,2406,2406,2406,2149,2149,1893,1876,1620,1347,1074,1074,818,802,818,1092,1638,1928,273,273,273,273,273},
'{273,273,273,273,273,273,273,2458,1895,1092,803,546,530,530,802,1075,1348,1621,1894,2150,2150,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2405,2149,2149,2149,2149,2149,2149,2149,2149,2405,2405,2405,2405,2388,2132,2132,2132,2132,2132,2132,2132,2132,2132,2116,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1586,1586,1586,1586,1586,1859,1859,2115,2132,2132,2132,2405,2405,2405,2405,2405,2405,2405,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2406,2149,2149,2149,2149,1876,1620,1347,1075,1074,802,802,802,1092,1382,1928,273,273,273,273,273},
'{273,273,273,273,273,273,273,2457,1639,1092,803,530,530,530,546,1075,1348,1621,1894,2150,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2133,2133,2133,2133,2133,2133,2133,2133,2405,2405,2405,2405,2404,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2116,2116,2116,2116,2116,2115,2115,2115,2115,2115,1859,1859,1859,1859,1843,1586,1586,1586,1586,1859,1859,2116,2132,2132,2132,2389,2405,2405,2405,2405,2405,2405,2405,2406,2405,2405,2405,2406,2406,2406,2406,2406,2406,2406,2422,2406,2405,2149,2149,2149,2149,1893,1876,1347,1331,1074,802,802,803,1092,1382,1912,273,273,273,273,273},
'{273,273,273,273,273,273,273,2457,1639,1092,803,530,530,530,802,1075,1348,1621,1894,2150,2149,2149,2149,2149,2133,2133,2133,2149,2133,2149,2149,2149,2133,2133,2133,2132,2132,2132,2132,2132,2132,2132,2132,2405,2405,2404,2388,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2116,2116,2115,2115,2115,2115,2115,2115,2115,2115,2115,2115,1859,1859,1859,1859,1859,1859,1859,1859,2116,2132,2132,2132,2132,2133,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2406,2406,2406,2406,2406,2406,2406,2406,2405,2149,2149,2149,2149,1893,1876,1604,1347,1074,802,802,802,1092,1382,1928,273,273,273,273,273},
'{273,273,273,273,273,273,273,2457,1639,1092,803,530,529,530,802,1075,1348,1621,1893,2150,2149,2149,2149,2133,2133,2132,2133,2133,2133,2133,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2404,2404,2388,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2116,2116,2115,2115,2115,2115,1843,1859,1859,1859,2115,2115,2115,2115,1859,1859,1859,1859,1859,2132,2132,2132,2132,2132,2133,2133,2133,2149,2149,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2406,2406,2406,2406,2149,2149,2149,2149,2149,1893,1877,1620,1347,1074,546,546,802,1092,1382,1928,273,273,273,273,273},
'{273,273,273,273,273,273,273,2457,1895,1092,819,546,529,546,802,1075,1348,1621,1893,1893,2149,2149,2149,2133,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2115,2115,1859,1859,1843,1843,1843,1843,1843,1843,1843,1843,1843,1843,1859,1859,1859,1859,1859,1859,1860,2116,2132,2132,2132,2132,2132,2389,2149,2149,2149,2149,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2149,2149,2405,2405,2149,2149,2149,2149,2149,2149,1877,1620,1347,1074,546,546,546,1092,1638,1928,273,273,273,273,273},
'{273,273,273,273,273,273,2971,2457,1895,1348,819,546,529,802,818,1075,1348,1621,1893,1893,2149,2149,2149,2149,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2116,2116,2115,1859,1859,1859,1842,1842,1842,1842,1842,1842,1842,1842,1842,1842,1842,1586,1842,1842,1843,1859,1859,2116,2132,2132,2132,2132,2132,2132,2132,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,1877,1620,1347,1074,545,546,546,1092,1638,2184,273,273,273,273,273},
'{273,273,273,273,273,273,2730,2441,1894,1348,1075,802,802,802,1075,1347,1620,1621,1877,1893,1893,2149,2149,2133,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2116,1859,1859,1859,1859,1859,1859,1843,1842,1586,1586,1570,1826,1826,1826,1826,1826,1826,1570,1570,1586,1586,1586,1842,1843,1859,1859,2116,2132,2132,2132,2132,2132,2132,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2405,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,2149,1877,1620,1347,1074,529,546,802,1092,1638,2185,273,273,273,273,273},
'{273,273,273,273,273,2730,2713,2440,1894,1604,1347,1074,1074,1075,1347,1348,1620,1877,1893,1893,2149,2149,2149,2149,2148,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1859,1859,1859,1859,1843,1842,1842,1586,1586,1586,1842,1842,1842,1843,1842,1842,1842,1842,1842,1586,1586,1586,1586,1842,1843,1859,1859,1859,1860,2132,2132,2132,2132,2133,2405,2405,2405,2405,2405,2405,2405,2405,2149,2133,2133,2132,2132,2148,2149,2149,2149,2149,2149,2149,2149,2149,2133,2149,2149,2149,1893,1877,1604,1347,1074,529,546,547,1092,1639,2185,273,273,273,273,273},
'{273,273,273,273,0,2713,2440,2167,1894,1620,1348,1347,1347,1347,1604,1620,1876,1877,1893,2149,2149,2133,2149,2132,2148,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1843,1586,1586,1586,1586,1842,1586,1586,1586,1586,1842,1842,1843,1843,0,0,0,0,0,0,0,0,0,0,1586,1586,1586,1843,1859,1859,1859,2132,2132,2132,2132,2133,2405,2405,2405,2405,2405,2405,2149,2133,2132,2132,2132,2132,2132,2132,2132,2133,2133,2133,2133,2133,2133,2133,2133,2149,2149,1877,1877,1604,1347,802,529,546,803,1092,1639,2185,273,273,273,273,273},
'{273,273,273,273,2696,2423,2151,2150,1877,1604,1603,1603,1603,1604,1620,1876,1876,1877,1877,2133,2133,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1859,1586,1586,1586,1586,1586,1586,1842,1842,1842,1842,1843,1843,0,0,0,0,0,0,0,0,0,0,0,0,0,1586,1586,1586,1587,1859,1859,1859,1860,2132,2132,2132,2133,2405,2405,2405,2405,2405,2149,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2133,2133,2133,2132,2132,2133,2133,1877,1877,1877,1604,1331,802,530,546,803,1093,1639,2185,273,273,273,273,273},
'{273,273,273,2696,2151,2133,1877,1860,1604,1603,1603,1876,1876,1876,1876,1876,1876,1877,2133,2133,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1586,1586,1586,1569,1570,1586,1586,1842,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1586,1587,1859,1859,1859,1859,2132,2132,2132,2132,2149,2149,2149,2405,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2133,1877,1877,1876,1604,1331,802,530,546,819,1093,1655,2186,273,273,273,273,273},
'{273,273,2696,2423,1877,1860,1603,1587,1587,1603,1603,1859,1860,1876,1876,1876,1876,1876,1877,1877,1877,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2131,1859,1859,1586,1586,1586,1586,1586,1586,1586,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1586,1586,1587,1603,1859,1859,1876,2132,2132,2149,2149,2149,2405,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1877,1877,1877,1620,1348,1331,802,530,546,819,1365,1911,2184,273,273,273,273,273},
'{273,2730,2423,2133,1860,1587,1570,1314,1586,1586,1603,1859,1859,1860,1876,1860,1860,1876,1876,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1859,1587,1586,1586,1586,1586,1843,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1586,1586,1586,1587,1859,1859,2132,2132,2132,2149,2149,2149,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1877,1877,1876,1604,1347,1075,802,530,803,820,1365,1912,0,273,273,273,273,273},
'{273,2423,2150,1860,1587,1570,1570,1570,1586,1586,1843,1859,1859,1859,1860,1860,1860,1876,1876,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1859,1859,1587,1843,1859,1859,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1314,1586,1586,1586,1603,1859,1876,2132,2132,2149,2149,2149,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1876,1876,1604,1331,1075,802,530,803,1076,1366,1912,273,273,273,273,273,273},
'{273,2423,1877,1859,1587,1586,1586,1586,1842,1842,1842,1859,1859,1859,1860,1860,1860,1876,1876,1876,1877,2132,2132,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1859,1859,1859,1859,1860,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1586,1586,1586,1587,1859,1860,2132,2132,2149,2149,2149,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1876,1876,1876,1604,1331,1058,802,530,819,1092,1638,2185,273,273,273,273,273,273},
'{273,2150,1860,1843,1842,1842,1842,1842,1842,1843,1843,1843,1859,1859,1860,1860,1860,1876,1876,1876,1877,2132,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1860,1860,1876,2132,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1586,1586,1586,1587,1859,1859,2132,2132,2132,2133,2149,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1876,1876,1604,1604,1331,1058,802,546,819,1349,1639,2185,273,273,273,273,273,273},
'{2184,2150,1860,1843,1842,1842,1842,2115,2115,2115,1859,1842,1859,1859,1860,1860,1860,1876,1876,1876,1876,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1587,1603,1603,1859,1859,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1876,1860,1604,1347,1075,1058,802,546,1076,1365,1911,2458,273,273,273,273,273,273},
'{2440,2150,1860,1843,1842,2098,2115,2115,2115,2115,1859,1842,1587,1859,1860,1860,1876,1620,1604,1876,1876,1876,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2131,2131,2132,2132,2132,2132,2132,2132,2132,2132,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1859,1859,1859,1859,1859,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,2132,1876,1876,1876,1876,1876,1860,1604,1331,1074,802,802,802,1076,1366,1912,2458,273,273,273,273,273,273},
'{2696,2406,1860,1843,1843,2099,2115,2115,2115,2115,1843,1586,1586,1603,1603,1860,1876,1876,1620,1876,1876,1876,1876,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,0,0,0,0,0,0,0,0,529,1041,1314,1586,1843,1843,1843,1842,1314,1057,528,0,0,0,0,0,0,0,0,0,0,1859,1859,1859,1860,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1876,1876,1876,1860,1604,1331,1074,1058,802,802,1348,1638,2184,2457,273,273,273,273,273,273},
'{2680,2406,2116,1859,2115,2115,2115,2116,2115,1859,1842,1586,1586,1603,1603,1603,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,0,0,0,256,529,1330,1586,1843,1843,2115,2115,2115,2115,2099,1843,1843,1843,1843,1843,1842,1314,785,0,0,0,0,0,0,0,0,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1876,1876,1876,1604,1604,1347,1330,1058,1058,1075,1349,1895,2441,3983,273,273,273,273,273,273},
'{2696,2406,2133,2116,2115,2115,2115,2116,2115,1843,1586,1330,1330,1586,1603,1603,1604,1620,1620,1876,1876,1876,1876,1876,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,0,0,529,1859,2132,1876,1859,2115,2115,2115,2115,2115,2115,2115,2115,2115,2115,2115,1859,1859,1859,1843,1586,785,256,0,0,0,0,0,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1860,1860,1876,1604,1604,1603,1331,1330,1331,1331,1621,1911,2440,2730,273,273,273,273,273,273},
'{2696,2406,2133,2116,2116,2115,2116,2116,1859,1842,1586,1313,1313,1330,1330,1603,1603,1604,1604,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1074,2132,2132,2132,2132,1859,1859,1859,1859,1843,1843,1843,1843,1843,1843,1843,1843,1843,1843,1843,1843,1586,1586,1586,1057,256,0,0,0,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1860,1860,1860,1860,1604,1604,1604,1603,1603,1603,1604,1877,2150,2440,2714,273,273,273,273,273,273},
'{2696,2422,2133,2132,2132,2115,2115,2115,1859,1586,1586,1313,1313,1330,1330,1587,1603,1604,1604,1860,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1843,1842,1842,1842,1842,1586,1842,1842,1842,1842,1843,1843,1843,1587,1586,1586,1586,1586,1330,529,0,0,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1860,1859,1603,1603,1603,1604,1604,1603,1603,1604,1604,1877,1894,2167,2440,273,273,273,273,273,273},
'{2696,2423,2405,2132,2132,2115,2115,2115,1842,1586,1313,1313,1313,1330,1330,1587,1603,1603,1860,1860,1860,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1876,1860,1860,1860,1860,2116,2132,2132,1876,1876,2132,2132,2132,2132,2132,2132,2133,2133,2133,2133,2133,2132,2132,2132,2132,1859,1843,1842,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1314,529,0,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1859,1859,1603,1603,1603,1603,1603,1603,1603,1604,1604,1876,1877,2150,2167,2440,273,273,273,273,273},
'{2696,2423,2405,2132,2132,2115,2115,1859,1842,1586,1569,1313,1313,1330,1586,1587,1603,1603,1860,1860,1860,1876,1876,1876,1876,1876,1876,1876,1876,1875,1859,1859,1859,1859,1859,1859,1860,1860,2116,2132,1876,1876,2132,2132,2132,2132,2132,2133,2149,2405,2405,2405,2405,2149,2133,2132,2132,1859,1586,1586,1586,1586,1586,1586,1586,1570,1570,1570,1570,1570,1570,1586,1586,1586,1586,1586,1586,1586,1314,1330,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1860,1859,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1604,1876,1894,2167,2440,273,273,273,273},
'{2696,2423,2149,2132,2132,2115,2115,1858,1842,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1860,1860,1860,1860,1860,1860,1860,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1860,1860,1860,2132,1876,1876,2132,2132,2132,2132,2132,2148,2149,2405,2405,2405,2405,2405,2149,2132,2132,1859,1587,1586,1586,1586,1586,1586,1586,1570,1570,1570,1570,1570,1570,1586,1586,1586,1586,1587,1586,1586,1586,1586,1859,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1860,1860,1859,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1603,1587,1603,1876,1894,2423,273,273,273,273},
'{2696,2422,2149,2132,2132,2115,2115,1842,1842,1842,1842,1859,1859,1859,1859,1859,1603,1603,1603,1603,1604,1860,1860,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1860,1860,2116,2132,2132,2132,2132,2132,2132,2148,2148,2149,2405,2405,2405,2405,2405,2149,2132,2132,1859,1859,1603,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1843,1843,1843,1859,1587,1587,1587,1859,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1860,1860,1860,1859,1859,1603,1603,1603,1603,1603,1603,1603,1858,1842,1586,1586,1586,1603,1876,2150,2730,273,273,273},
'{2440,2423,2149,2132,2132,2115,2115,2115,2115,1859,2115,2115,2115,2115,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1860,1860,1876,2132,2132,2132,2132,2132,2132,2148,2149,2149,2405,2405,2405,2405,2405,2149,2132,2132,1859,1859,1859,1859,1859,1587,1587,1586,1586,1586,1586,1586,1587,1843,1843,1859,1859,1859,1859,1859,1859,1859,1859,1859,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1860,1860,1860,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1858,1858,1842,1586,1586,1587,1860,2150,2440,273,273,273},
'{2184,2423,2149,2132,2132,2115,2115,2115,2115,2115,2132,2388,2132,2132,2132,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1860,1860,1876,2132,2132,2132,2132,2132,2132,2132,2149,2149,2405,2405,2405,2405,2405,2149,2132,2132,1876,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1860,1860,1860,1859,1876,2132,2132,2132,2132,2132,2132,2132,1876,2132,2132,2132,2132,1876,1876,1876,1876,1876,1860,1860,1859,1859,1859,1603,1603,1603,1603,1603,1602,1602,1602,1603,1859,2114,1842,1842,1586,1587,1860,2150,2440,273,273,273},
'{273,2439,2150,2133,2132,2116,2115,2115,2116,2132,2132,2388,2132,2132,2132,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1860,1860,1876,2132,2132,2132,2132,2132,2132,2132,2132,2149,2149,2149,2405,2405,2149,2132,2132,2132,1876,1876,1860,1860,1876,1876,2132,1876,1860,1859,1859,1859,1859,1859,1859,1859,1859,1860,2116,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1876,1876,1876,1876,1876,1876,1860,1860,1860,1876,1860,1860,1859,1859,1603,1603,1603,1603,1587,1586,1586,1602,1603,1859,1859,2115,1859,1842,1843,1859,1860,2150,2424,273,273,273},
'{273,2440,2166,2149,2132,2116,2116,2116,2132,2132,2132,2132,2132,2115,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1860,1860,1860,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2149,2149,2149,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1860,1860,1860,1860,1860,2116,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2131,1875,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1586,1586,1586,1586,1602,1603,1859,1859,2115,2115,1859,1859,1859,1860,2150,2424,273,273,273},
'{273,2184,2423,2150,2133,2132,2132,2132,2132,2132,2132,2116,1859,1859,1859,1603,1586,1586,1330,1347,1347,1347,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1860,1860,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2131,1875,1875,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1587,1586,1330,1586,1586,1586,1859,1859,2115,2115,2115,2115,1859,1860,1860,2150,2440,273,273,273},
'{273,273,2697,2423,2150,2133,2133,1876,1876,1860,1860,1859,1859,1587,1587,1586,1330,1330,1330,1330,1330,1331,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1876,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2131,1875,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1587,1586,1330,1330,1330,1586,1586,1603,1859,1859,2115,2116,2116,2116,1860,2133,2407,2696,273,273,273},
'{273,273,273,2440,2167,2150,2133,1877,1876,1860,1860,1603,1587,1587,1330,1330,1314,1330,1330,1330,1330,1330,1347,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1860,1876,1876,1876,1876,1876,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2131,1875,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1587,1586,1330,1330,1330,1330,1586,1603,1859,1859,2116,2116,2116,2116,2116,2133,2423,2697,273,273,273},
'{273,273,273,273,2440,2423,2167,2150,1877,1877,1860,1604,1603,1587,1587,1330,1314,1314,1058,1330,1330,1331,1331,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,2133,2149,2133,2133,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1875,1875,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1587,1587,1586,1330,1314,1314,1314,1330,1587,1859,1859,2116,2116,2116,2116,2133,2134,2424,2713,273,273,273},
'{273,273,273,273,273,2457,2440,2167,1894,1877,1877,1860,1604,1603,1587,1330,1314,1314,1058,1330,1331,1331,1331,1587,1587,1587,1587,1603,1603,1603,1586,1586,1586,1586,1586,1587,1587,1587,1587,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,2405,2405,2405,2149,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1858,1858,1858,1602,1586,1586,1586,1587,1587,1587,1587,1330,1314,1314,1314,1330,1586,1603,1859,2116,2116,2116,2117,2133,2406,2440,273,273,273,273},
'{273,273,273,273,273,273,273,2440,2168,2167,1894,1894,1878,1877,1877,1348,1074,1058,1058,1074,1331,1331,1331,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1587,1587,1587,1587,1603,1603,1603,1603,1603,1603,1603,1859,2405,2405,2405,2149,2148,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1858,1858,1602,1602,1858,1858,1602,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1586,1586,1603,1859,2116,2116,2116,2133,2134,2407,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,2184,2184,2167,2167,1911,1621,1075,1075,1058,1074,1331,1331,1331,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1587,1587,1587,1587,1587,1587,1587,1587,1587,1859,2405,2405,2405,2149,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1876,1859,1859,1859,1859,1859,1859,1859,1859,1858,1858,1586,1586,1586,1586,1858,1858,1586,1586,1586,1586,1586,1586,1330,1330,1330,1586,1587,1586,1586,1586,1586,1842,1859,2115,2116,2116,2133,2406,2440,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1638,1076,1075,1074,1074,1331,1331,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1587,1587,1587,1587,1587,1587,1330,1603,2405,2405,2405,2405,2132,2132,2132,2132,2132,2132,2132,1860,1859,1859,1859,2131,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1603,1603,1603,1859,1859,1859,1859,1859,1602,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1586,1587,1587,1587,1842,1842,1843,1859,2115,2116,2116,2133,2406,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1894,1348,1075,1075,1075,1331,1331,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,2149,2405,2149,2132,2132,2132,2132,2132,2132,1876,1860,1859,1859,1859,1859,1859,1875,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,2132,1859,1586,1586,1586,1587,1603,1603,1603,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1586,1587,1859,1859,1859,1859,1859,2115,2116,2116,2132,2149,2423,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1365,1092,1075,1075,1075,1331,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1586,2132,2132,2132,2132,2132,2132,1876,1876,1860,1859,1859,1859,1859,1859,1859,1859,1859,1876,2132,2132,2132,2132,2132,2132,2132,2132,1859,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1586,1586,1859,1859,1859,2115,2115,2116,2116,2132,2133,2150,2423,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1638,1349,1075,1075,1075,1075,1331,1331,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1330,1330,1330,1314,1314,1314,1314,1314,1314,1314,1603,2132,2132,1876,1876,1860,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1860,1876,2132,2132,2132,2132,2132,2132,2132,1586,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1587,1859,1859,2115,2115,2116,2116,2133,2133,2150,2184,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1895,1365,1075,1075,1075,1075,1331,1347,1331,1330,1330,1330,1330,1330,1330,1330,1330,1074,1074,1074,1058,1058,1058,1314,1314,1314,1314,1314,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1330,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1860,2132,2132,2132,2132,2132,2132,1586,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1330,1330,1330,1586,1586,1330,1330,1330,1330,1330,1330,1330,1074,1058,1058,1058,1330,1330,1330,1330,1586,1859,1859,2115,2132,2132,1860,1877,2133,2150,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1638,1092,1075,1075,1075,1331,1347,1331,1331,1331,1330,1330,1330,1330,1074,1074,1074,1074,1074,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1314,1314,1330,1586,1587,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1860,2132,2132,2132,1876,1330,1314,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1074,1058,1058,1074,1331,1331,1603,1603,1603,1603,1859,1859,1860,1860,1876,1877,2150,2184,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1639,1349,1092,1076,1075,1347,1347,1331,1331,1331,1330,1330,1074,1074,1074,1074,1074,1074,1058,1058,1058,1058,1058,1058,1074,1074,1074,1074,1074,1074,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1314,1314,1314,1314,1314,1314,1314,1330,1330,1330,1586,1586,1587,1587,1603,1603,1603,1587,1058,1058,1058,1058,1314,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1074,1058,1058,1058,1075,1331,1604,1604,1877,1604,1603,1587,1603,1860,1860,1877,1877,2150,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1911,1365,1348,1348,1348,1347,1347,1347,1331,1331,1331,1330,1074,1074,1074,1074,1074,1074,1074,1058,1058,1058,1058,1058,1074,1074,1074,1074,1074,1074,1074,1074,1058,1058,1058,1058,1058,1058,1058,1058,1314,1314,1314,1314,1314,1314,1314,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1074,1074,1074,1074,1075,1075,1348,1894,1894,2150,1894,1621,1604,1604,1860,1877,1894,2150,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1638,1365,1348,1348,1348,1347,1347,1331,1331,1331,1331,1331,1074,1074,1074,1074,1074,1074,1058,1058,1058,1058,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1058,1058,1058,1058,1058,1058,1058,1314,1314,1314,1314,1314,1314,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1074,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1074,1074,1075,1075,1075,1348,1622,2167,2440,2184,2168,1894,1878,1877,1877,1894,2167,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1895,1622,1349,1348,1348,1347,1347,1331,1331,1331,1331,1331,1331,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1058,1058,1058,1058,1058,1058,1314,1314,1314,1314,1314,1314,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1074,1330,1330,1330,1330,1074,1074,1074,1074,1074,1074,1074,1074,1074,1330,1074,1075,1075,1075,1075,1092,1365,1911,2184,273,273,273,273,2184,1895,1895,4095,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1641,1894,1621,1348,1348,1348,1347,1347,1331,1331,1331,1331,1331,1330,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1074,1330,1074,1074,1074,1074,1074,1058,1058,1058,1058,1058,1314,1314,1314,1314,1314,1314,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1074,1074,1074,1075,1075,1075,1076,1349,1638,2457,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1911,1622,1349,1348,1348,1347,1347,1331,1331,1331,1331,1331,1330,1330,1330,1330,1074,1074,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1058,1058,1058,1314,1314,1314,1314,1314,1314,1314,1314,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1074,1074,1075,1075,1075,1092,1366,1912,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2168,1894,1621,1620,1604,1604,1603,1347,1331,1331,1331,1331,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1074,1075,1075,1092,1366,1911,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1895,1622,1621,1604,1604,1603,1603,1587,1331,1331,1331,1331,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1330,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1075,1092,1365,1639,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2168,1894,1877,1604,1604,1603,1603,1587,1587,1587,1331,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1330,1330,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1075,1075,1348,1638,2184,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1895,1877,1620,1604,1604,1603,1587,1587,1587,1587,1587,1587,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1314,1058,1058,1314,1314,1314,1314,1314,1314,1314,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1074,1075,1075,1075,1076,1365,1911,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2440,2167,1893,1876,1604,1604,1603,1603,1587,1587,1587,1587,1587,1587,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1330,1330,1330,1330,1314,1330,1330,1330,1330,1330,1330,1330,1314,1330,1074,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1058,1074,1075,1075,1348,1348,1638,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2440,2167,1894,1876,1876,1604,1604,1603,1603,1603,1587,1587,1587,1587,1587,1587,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1330,1314,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1330,1074,1058,1058,1058,1058,1058,1058,1058,1058,1058,1074,1330,1075,1331,1348,1621,2409,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2730,2167,2150,1876,1876,1860,1604,1603,1603,1603,1603,1587,1587,1587,1587,1587,1331,1331,1331,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1314,1314,1314,1058,1058,1058,1314,1314,1314,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1058,1058,1058,1058,1058,1074,1330,1330,1330,1331,1331,1621,1894,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,2167,2150,1876,1876,1860,1604,1603,1603,1603,1603,1587,1587,1587,1587,1587,1587,1587,1331,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1314,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1074,1074,1074,1058,1074,1074,1330,1330,1331,1331,1348,1621,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,2150,1876,1876,1860,1604,1604,1603,1603,1603,1603,1587,1587,1587,1587,1587,1587,1587,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1314,1314,1314,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1074,1074,1074,1074,1330,1330,1331,1331,1347,1348,1622,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,2150,1876,1876,1860,1604,1603,1603,1603,1603,1603,1587,1587,1587,1587,1587,1587,1587,1587,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1314,1314,1314,1314,1314,1314,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1074,1074,1074,1074,1330,1330,1331,1331,1331,1347,1604,1894,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,2150,1876,1876,1860,1860,1603,1603,1603,1603,1603,1587,1587,1587,1587,1587,1587,1587,1587,1587,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1331,1331,1331,1347,1348,1620,1894,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,2150,1876,1876,1876,1860,1603,1603,1603,1603,1603,1603,1603,1587,1587,1587,1587,1587,1587,1587,1587,1587,1331,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1331,1331,1331,1331,1347,1604,1621,1894,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,2149,1876,1876,1876,1860,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1587,1587,1587,1587,1587,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1331,1331,1331,1347,1603,1604,1621,1894,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,2149,1876,1876,1876,1860,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1587,1587,1587,1587,1587,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1331,1331,1331,1603,1603,1604,1621,1894,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,1893,1876,1876,1876,1860,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1587,1587,1587,1587,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1587,1603,1603,1603,1604,1621,1894,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,1893,1876,1876,1876,1860,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1587,1587,1587,1587,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1603,1603,1603,1603,1620,1621,1911,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2166,1893,1876,1876,1876,1860,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1587,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1620,1621,1911,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,0,2166,1893,1876,1876,1876,1860,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1602,1603,1603,1603,1603,1603,1620,1621,1911,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,4095,2166,1893,1876,1876,1876,1876,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1620,1621,1911,0,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2730,2150,1893,1876,1876,1876,1876,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1859,1603,1620,1637,1911,4095,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2457,2150,1893,1876,1876,1876,1876,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1603,1859,1603,1620,1637,1911,4095,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,2150,1893,1876,1876,1876,1876,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1587,1587,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1604,1620,1894,1911,2184,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,1894,1893,1876,1876,1876,1876,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1587,1603,1587,1587,1587,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1620,1620,1637,1911,1365,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,1894,1893,1876,1876,1876,1876,1859,1859,1859,1859,1859,1603,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1876,1620,1637,1911,2730,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,1894,1877,1876,1876,1876,1860,1859,1859,1859,1859,1859,1603,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1876,1620,1637,1911,1638,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2167,1894,1877,1876,1876,1876,1860,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1876,1876,1893,1910,2406,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1911,1894,1877,1876,1876,1876,1860,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1876,1876,1893,1910,2184,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1911,1894,1877,1876,1876,1876,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1876,1876,1893,1910,2167,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,1911,1894,1877,1876,1876,1876,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1876,1876,1893,1894,2184,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,2184,2167,1911,1894,1877,1876,1876,1860,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1876,1876,1877,1894,2168,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1912,1911,1911,1894,1894,1877,1876,1876,1860,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1876,1876,1877,1894,2168,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1656,1639,1639,1638,1894,1893,1877,1876,1876,1860,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1876,1876,1621,1894,2168,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,273},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,273,1384,1367,1366,1366,1622,1621,1877,1876,1876,1876,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1876,1876,1621,1895,1912,273,273,273,273,273,273,273,273,273,2184,1657,1657,1657,1657,1657,1657,1641,1641,1384,1384,1385,1385,1641,1657,1657,1658},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,273,1384,1111,1093,1093,1093,1349,1621,1621,1876,1876,1876,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1876,1877,1621,1895,1912,1641,273,273,273,273,273,273,1657,1401,1385,1384,1384,1385,1385,1384,1384,1368,1368,1112,1112,1112,1112,1384,1385,1657,1658},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,1657,1111,1094,821,821,1092,1348,1621,1621,1876,1876,1876,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1860,1620,1621,1894,1896,1913,273,273,273,273,1675,1674,1402,1385,1385,1129,1112,1113,1113,1368,1368,1112,1112,1095,1095,1095,1112,1112,1385,1657,1658},
'{273,273,273,273,273,273,273,273,273,273,273,273,273,1384,1094,821,548,820,1076,1348,1605,1620,1876,1876,1876,1859,1859,1875,1875,1875,1875,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1586,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1876,1620,1621,1622,1895,1912,1913,1930,1674,1675,1675,1659,1402,1385,1129,1113,1112,1113,1113,1112,1112,1096,839,839,839,839,839,1112,1385,1401,1658},
'{273,273,273,273,273,273,273,273,273,273,273,273,1913,1368,838,821,548,820,1076,1348,1604,1876,1876,1876,1876,1859,1859,1875,1875,1875,1875,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1860,1604,1621,1622,1639,1640,1657,1658,1658,1659,1659,1659,1402,1386,1385,1113,1113,1113,1113,1112,1112,840,839,839,839,839,840,1112,1385,1658,1931},
'{273,273,273,273,273,273,273,273,273,273,273,273,1657,1111,821,821,548,820,1348,1604,1620,1876,1876,1876,1876,1859,1859,1859,1859,1875,1875,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1587,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1587,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1604,1604,1621,1622,1639,1640,1641,1658,1658,1659,1659,1402,1402,1386,1129,1113,1113,1113,1112,1112,856,840,839,839,839,856,1113,1386,1658,1931},
'{273,273,273,273,273,273,273,273,273,273,273,4095,1640,1095,821,548,547,820,1348,1604,1876,1876,1876,1876,1876,1859,1859,1859,1859,1875,1875,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1587,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1604,1604,1621,1622,1623,1640,1641,1641,1658,1658,1659,1402,1402,1386,1129,1113,1113,1113,1113,1112,856,840,840,840,840,1112,1113,1402,1931,1948},
'{273,273,273,273,273,273,273,273,273,273,273,1914,1384,1094,549,548,547,1076,1348,1604,1876,1876,1876,1876,1875,1859,1859,1859,1859,1875,1875,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1876,1876,1876,1876,1859,1859,1859,1859,1859,1859,1604,1620,1621,1622,1367,1384,1385,1386,1402,1658,1402,1402,1386,1129,1113,1113,1113,1113,1113,857,856,840,840,840,1113,1385,1658,1931,2204},
'{273,273,273,273,273,273,273,273,273,273,273,1657,1367,822,548,548,547,1076,1348,1604,1876,1876,1876,1876,1875,1859,1859,1859,1859,1875,1875,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1330,1330,1330,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1876,1876,1876,1876,1876,1859,1859,1859,1859,1859,1859,1860,1620,1621,1622,1367,1367,1384,1385,1401,1658,1402,1386,1385,1113,1113,1113,1113,1113,1113,1113,857,856,856,856,1113,1386,1659,1932,2204},
'{273,273,273,273,273,273,273,273,273,273,273,1640,1367,821,548,804,803,1076,1604,1604,1876,1876,1876,1876,1875,1875,1875,1875,1875,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1586,1586,1586,1586,1586,1330,1330,1330,1330,1330,1586,1586,1586,1586,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1876,1876,1876,1876,1876,1876,1875,1859,1859,1859,1859,1859,1860,1604,1621,1621,1622,1623,1639,1640,1641,1641,1641,1385,1385,1113,1112,1112,1112,1113,1113,1113,856,856,856,1113,1385,1658,1931,2204,2204},
'{273,273,273,273,273,273,273,273,273,273,2184,1384,1094,820,803,803,1076,1348,1604,1876,1876,1876,1876,1876,1876,1876,1875,1875,1875,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1586,1586,1586,1586,1586,1586,1330,1330,1330,1330,1586,1586,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1875,1876,1876,1876,1876,1876,1876,1876,1876,1859,1859,1859,1859,1859,1860,1860,1604,1621,1621,1622,1623,1623,1640,1640,1640,1624,1368,1368,1112,1112,1112,1112,1112,1112,856,1112,1113,1129,1386,1658,1931,2204,2204},
'{273,273,273,273,273,273,273,273,273,273,1929,1383,1094,820,803,1075,1332,1604,1604,1876,1876,1876,1876,1876,1876,1876,1875,1875,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1875,1876,1876,1876,1876,1876,1876,1876,1876,1859,1859,1859,1859,1859,1859,1860,1860,1621,1621,1622,1878,1879,1623,1623,1623,1368,1368,1367,1095,1095,839,840,1096,1096,840,1112,1113,1385,1402,1675,1931,2204,2204},
'{273,273,273,273,273,273,273,273,273,273,1657,1383,1094,1076,803,1075,1348,1604,1876,1876,1876,1876,1876,1875,1875,1875,1875,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1875,1876,1876,1876,1876,1876,1876,1876,1876,1859,1859,1859,1859,1859,1859,1859,1860,1860,1877,1877,1878,1878,1622,1623,1623,1367,1351,1095,1095,839,823,839,839,840,840,1096,1112,1385,1658,1931,1932,2204,2220},
'{273,273,273,273,273,273,273,273,273,273,1657,1367,1093,1076,1075,1331,1604,1604,1876,1876,1876,1876,1876,1875,1875,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1587,1586,1586,1586,1586,1586,1586,1586,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1875,1876,1876,1876,1876,1876,1876,1876,1876,1859,1859,1859,1859,1859,1859,1859,1860,1860,1876,1877,1877,1877,1878,1622,1622,1606,1350,1094,1094,822,822,822,839,839,839,1096,1112,1385,1658,1931,1948,2204,2220},
'{273,273,273,273,273,273,273,273,273,273,1657,1367,1093,1076,1075,1347,1604,1876,1876,1876,1876,1876,1876,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1859,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1587,1586,1586,1586,1586,1586,1586,1586,1586,1587,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1603,1859,1859,1859,1859,1859,1859,1859,1875,1876,1876,1876,1876,1876,1876,1876,1876,1859,1859,1859,1859,1859,1859,1859,1859,1860,1876,1876,1877,1877,1877,1877,1621,1605,1349,1349,1077,1077,821,822,822,823,1095,1096,1368,1385,1658,1931,1948,2204,2204}
};



endmodule